// Generator : SpinalHDL v1.7.2    git head : 08fc866bebdc40c471ebe327bface63e34406489
// Component : SystolicArray
// Date      : 09/12/2022, 23:09:14

`timescale 1ns/1ps

module SystolicArray (
  input               start,
  input               last,
  input      [511:0]  A_Array,
  input      [511:0]  B_Array,
  output reg [2047:0] Array_OUT,
  input               clk,
  input               reset
);

  wire       [63:0]   tile_8_A;
  wire       [63:0]   tile_8_B;
  wire       [63:0]   tile_9_A;
  wire       [63:0]   tile_9_B;
  wire       [63:0]   tile_10_A;
  wire       [63:0]   tile_10_B;
  wire       [63:0]   tile_11_A;
  wire       [63:0]   tile_11_B;
  wire       [63:0]   tile_12_A;
  wire       [63:0]   tile_12_B;
  wire       [63:0]   tile_13_A;
  wire       [63:0]   tile_13_B;
  wire       [63:0]   tile_14_A;
  wire       [63:0]   tile_14_B;
  wire       [63:0]   tile_15_A;
  wire       [63:0]   tile_15_B;
  wire       [2047:0] tile_8_Tile_OUT;
  wire       [2047:0] tile_9_Tile_OUT;
  wire       [2047:0] tile_10_Tile_OUT;
  wire       [2047:0] tile_11_Tile_OUT;
  wire       [2047:0] tile_12_Tile_OUT;
  wire       [2047:0] tile_13_Tile_OUT;
  wire       [2047:0] tile_14_Tile_OUT;
  wire       [2047:0] tile_15_Tile_OUT;
  wire       [31:0]   _zz_Array_OUT;
  wire       [31:0]   _zz_Array_OUT_1;
  wire       [31:0]   _zz_Array_OUT_2;
  wire       [31:0]   _zz_Array_OUT_3;
  wire       [31:0]   _zz_Array_OUT_4;
  wire       [31:0]   _zz_Array_OUT_5;
  wire       [31:0]   _zz_Array_OUT_6;
  wire       [31:0]   _zz_Array_OUT_7;
  wire       [31:0]   _zz_Array_OUT_8;
  wire       [31:0]   _zz_Array_OUT_9;
  wire       [31:0]   _zz_Array_OUT_10;
  wire       [31:0]   _zz_Array_OUT_11;
  wire       [31:0]   _zz_Array_OUT_12;
  wire       [31:0]   _zz_Array_OUT_13;
  wire       [31:0]   _zz_Array_OUT_14;
  wire       [31:0]   _zz_Array_OUT_15;
  wire       [31:0]   _zz_Array_OUT_16;
  wire       [31:0]   _zz_Array_OUT_17;
  wire       [31:0]   _zz_Array_OUT_18;
  wire       [31:0]   _zz_Array_OUT_19;
  wire       [31:0]   _zz_Array_OUT_20;
  wire       [31:0]   _zz_Array_OUT_21;
  wire       [31:0]   _zz_Array_OUT_22;
  wire       [31:0]   _zz_Array_OUT_23;
  wire       [31:0]   _zz_Array_OUT_24;
  wire       [31:0]   _zz_Array_OUT_25;
  wire       [31:0]   _zz_Array_OUT_26;
  wire       [31:0]   _zz_Array_OUT_27;
  wire       [31:0]   _zz_Array_OUT_28;
  wire       [31:0]   _zz_Array_OUT_29;
  wire       [31:0]   _zz_Array_OUT_30;
  wire       [31:0]   _zz_Array_OUT_31;
  wire       [31:0]   _zz_Array_OUT_32;
  wire       [31:0]   _zz_Array_OUT_33;
  wire       [31:0]   _zz_Array_OUT_34;
  wire       [31:0]   _zz_Array_OUT_35;
  wire       [31:0]   _zz_Array_OUT_36;
  wire       [31:0]   _zz_Array_OUT_37;
  wire       [31:0]   _zz_Array_OUT_38;
  wire       [31:0]   _zz_Array_OUT_39;
  wire       [31:0]   _zz_Array_OUT_40;
  wire       [31:0]   _zz_Array_OUT_41;
  wire       [31:0]   _zz_Array_OUT_42;
  wire       [31:0]   _zz_Array_OUT_43;
  wire       [31:0]   _zz_Array_OUT_44;
  wire       [31:0]   _zz_Array_OUT_45;
  wire       [31:0]   _zz_Array_OUT_46;
  wire       [31:0]   _zz_Array_OUT_47;
  wire       [31:0]   _zz_Array_OUT_48;
  wire       [31:0]   _zz_Array_OUT_49;
  wire       [31:0]   _zz_Array_OUT_50;
  wire       [31:0]   _zz_Array_OUT_51;
  wire       [31:0]   _zz_Array_OUT_52;
  wire       [31:0]   _zz_Array_OUT_53;
  wire       [31:0]   _zz_Array_OUT_54;
  wire       [31:0]   _zz_Array_OUT_55;
  wire       [31:0]   _zz_Array_OUT_56;
  wire       [31:0]   _zz_Array_OUT_57;
  wire       [31:0]   _zz_Array_OUT_58;
  wire       [31:0]   _zz_Array_OUT_59;
  wire       [31:0]   _zz_Array_OUT_60;
  wire       [31:0]   _zz_Array_OUT_61;
  wire       [31:0]   _zz_Array_OUT_62;
  wire       [31:0]   _zz_Array_OUT_63;
  wire       [31:0]   _zz_Array_OUT_64;
  wire       [31:0]   _zz_Array_OUT_65;
  wire       [31:0]   _zz_Array_OUT_66;
  wire       [31:0]   _zz_Array_OUT_67;
  wire       [31:0]   _zz_Array_OUT_68;
  wire       [31:0]   _zz_Array_OUT_69;
  wire       [31:0]   _zz_Array_OUT_70;
  wire       [31:0]   _zz_Array_OUT_71;
  wire       [31:0]   _zz_Array_OUT_72;
  wire       [31:0]   _zz_Array_OUT_73;
  wire       [31:0]   _zz_Array_OUT_74;
  wire       [31:0]   _zz_Array_OUT_75;
  wire       [31:0]   _zz_Array_OUT_76;
  wire       [31:0]   _zz_Array_OUT_77;
  wire       [31:0]   _zz_Array_OUT_78;
  wire       [31:0]   _zz_Array_OUT_79;
  wire       [31:0]   _zz_Array_OUT_80;
  wire       [31:0]   _zz_Array_OUT_81;
  wire       [31:0]   _zz_Array_OUT_82;
  wire       [31:0]   _zz_Array_OUT_83;
  wire       [31:0]   _zz_Array_OUT_84;
  wire       [31:0]   _zz_Array_OUT_85;
  wire       [31:0]   _zz_Array_OUT_86;
  wire       [31:0]   _zz_Array_OUT_87;
  wire       [31:0]   _zz_Array_OUT_88;
  wire       [31:0]   _zz_Array_OUT_89;
  wire       [31:0]   _zz_Array_OUT_90;
  wire       [31:0]   _zz_Array_OUT_91;
  wire       [31:0]   _zz_Array_OUT_92;
  wire       [31:0]   _zz_Array_OUT_93;
  wire       [31:0]   _zz_Array_OUT_94;
  wire       [31:0]   _zz_Array_OUT_95;
  wire       [31:0]   _zz_Array_OUT_96;
  wire       [31:0]   _zz_Array_OUT_97;
  wire       [31:0]   _zz_Array_OUT_98;
  wire       [31:0]   _zz_Array_OUT_99;
  wire       [31:0]   _zz_Array_OUT_100;
  wire       [31:0]   _zz_Array_OUT_101;
  wire       [31:0]   _zz_Array_OUT_102;
  wire       [31:0]   _zz_Array_OUT_103;
  wire       [31:0]   _zz_Array_OUT_104;
  wire       [31:0]   _zz_Array_OUT_105;
  wire       [31:0]   _zz_Array_OUT_106;
  wire       [31:0]   _zz_Array_OUT_107;
  wire       [31:0]   _zz_Array_OUT_108;
  wire       [31:0]   _zz_Array_OUT_109;
  wire       [31:0]   _zz_Array_OUT_110;
  wire       [31:0]   _zz_Array_OUT_111;
  wire       [31:0]   _zz_Array_OUT_112;
  wire       [31:0]   _zz_Array_OUT_113;
  wire       [31:0]   _zz_Array_OUT_114;
  wire       [31:0]   _zz_Array_OUT_115;
  wire       [31:0]   _zz_Array_OUT_116;
  wire       [31:0]   _zz_Array_OUT_117;
  wire       [31:0]   _zz_Array_OUT_118;
  wire       [31:0]   _zz_Array_OUT_119;
  wire       [31:0]   _zz_Array_OUT_120;
  wire       [31:0]   _zz_Array_OUT_121;
  wire       [31:0]   _zz_Array_OUT_122;
  wire       [31:0]   _zz_Array_OUT_123;
  wire       [31:0]   _zz_Array_OUT_124;
  wire       [31:0]   _zz_Array_OUT_125;
  wire       [31:0]   _zz_Array_OUT_126;
  wire       [31:0]   _zz_Array_OUT_127;
  wire       [31:0]   _zz_Array_OUT_128;
  wire       [31:0]   _zz_Array_OUT_129;
  wire       [31:0]   _zz_Array_OUT_130;
  wire       [31:0]   _zz_Array_OUT_131;
  wire       [31:0]   _zz_Array_OUT_132;
  wire       [31:0]   _zz_Array_OUT_133;
  wire       [31:0]   _zz_Array_OUT_134;
  wire       [31:0]   _zz_Array_OUT_135;
  wire       [31:0]   _zz_Array_OUT_136;
  wire       [31:0]   _zz_Array_OUT_137;
  wire       [31:0]   _zz_Array_OUT_138;
  wire       [31:0]   _zz_Array_OUT_139;
  wire       [31:0]   _zz_Array_OUT_140;
  wire       [31:0]   _zz_Array_OUT_141;
  wire       [31:0]   _zz_Array_OUT_142;
  wire       [31:0]   _zz_Array_OUT_143;
  wire       [31:0]   _zz_Array_OUT_144;
  wire       [31:0]   _zz_Array_OUT_145;
  wire       [31:0]   _zz_Array_OUT_146;
  wire       [31:0]   _zz_Array_OUT_147;
  wire       [31:0]   _zz_Array_OUT_148;
  wire       [31:0]   _zz_Array_OUT_149;
  wire       [31:0]   _zz_Array_OUT_150;
  wire       [31:0]   _zz_Array_OUT_151;
  wire       [31:0]   _zz_Array_OUT_152;
  wire       [31:0]   _zz_Array_OUT_153;
  wire       [31:0]   _zz_Array_OUT_154;
  wire       [31:0]   _zz_Array_OUT_155;
  wire       [31:0]   _zz_Array_OUT_156;
  wire       [31:0]   _zz_Array_OUT_157;
  wire       [31:0]   _zz_Array_OUT_158;
  wire       [31:0]   _zz_Array_OUT_159;
  wire       [31:0]   _zz_Array_OUT_160;
  wire       [31:0]   _zz_Array_OUT_161;
  wire       [31:0]   _zz_Array_OUT_162;
  wire       [31:0]   _zz_Array_OUT_163;
  wire       [31:0]   _zz_Array_OUT_164;
  wire       [31:0]   _zz_Array_OUT_165;
  wire       [31:0]   _zz_Array_OUT_166;
  wire       [31:0]   _zz_Array_OUT_167;
  wire       [31:0]   _zz_Array_OUT_168;
  wire       [31:0]   _zz_Array_OUT_169;
  wire       [31:0]   _zz_Array_OUT_170;
  wire       [31:0]   _zz_Array_OUT_171;
  wire       [31:0]   _zz_Array_OUT_172;
  wire       [31:0]   _zz_Array_OUT_173;
  wire       [31:0]   _zz_Array_OUT_174;
  wire       [31:0]   _zz_Array_OUT_175;
  wire       [31:0]   _zz_Array_OUT_176;
  wire       [31:0]   _zz_Array_OUT_177;
  wire       [31:0]   _zz_Array_OUT_178;
  wire       [31:0]   _zz_Array_OUT_179;
  wire       [31:0]   _zz_Array_OUT_180;
  wire       [31:0]   _zz_Array_OUT_181;
  wire       [31:0]   _zz_Array_OUT_182;
  wire       [31:0]   _zz_Array_OUT_183;
  wire       [31:0]   _zz_Array_OUT_184;
  wire       [31:0]   _zz_Array_OUT_185;
  wire       [31:0]   _zz_Array_OUT_186;
  wire       [31:0]   _zz_Array_OUT_187;
  wire       [31:0]   _zz_Array_OUT_188;
  wire       [31:0]   _zz_Array_OUT_189;
  wire       [31:0]   _zz_Array_OUT_190;
  wire       [31:0]   _zz_Array_OUT_191;
  wire       [31:0]   _zz_Array_OUT_192;
  wire       [31:0]   _zz_Array_OUT_193;
  wire       [31:0]   _zz_Array_OUT_194;
  wire       [31:0]   _zz_Array_OUT_195;
  wire       [31:0]   _zz_Array_OUT_196;
  wire       [31:0]   _zz_Array_OUT_197;
  wire       [31:0]   _zz_Array_OUT_198;
  wire       [31:0]   _zz_Array_OUT_199;
  wire       [31:0]   _zz_Array_OUT_200;
  wire       [31:0]   _zz_Array_OUT_201;
  wire       [31:0]   _zz_Array_OUT_202;
  wire       [31:0]   _zz_Array_OUT_203;
  wire       [31:0]   _zz_Array_OUT_204;
  wire       [31:0]   _zz_Array_OUT_205;
  wire       [31:0]   _zz_Array_OUT_206;
  wire       [31:0]   _zz_Array_OUT_207;
  wire       [31:0]   _zz_Array_OUT_208;
  wire       [31:0]   _zz_Array_OUT_209;
  wire       [31:0]   _zz_Array_OUT_210;
  wire       [31:0]   _zz_Array_OUT_211;
  wire       [31:0]   _zz_Array_OUT_212;
  wire       [31:0]   _zz_Array_OUT_213;
  wire       [31:0]   _zz_Array_OUT_214;
  wire       [31:0]   _zz_Array_OUT_215;
  wire       [31:0]   _zz_Array_OUT_216;
  wire       [31:0]   _zz_Array_OUT_217;
  wire       [31:0]   _zz_Array_OUT_218;
  wire       [31:0]   _zz_Array_OUT_219;
  wire       [31:0]   _zz_Array_OUT_220;
  wire       [31:0]   _zz_Array_OUT_221;
  wire       [31:0]   _zz_Array_OUT_222;
  wire       [31:0]   _zz_Array_OUT_223;
  wire       [31:0]   _zz_Array_OUT_224;
  wire       [31:0]   _zz_Array_OUT_225;
  wire       [31:0]   _zz_Array_OUT_226;
  wire       [31:0]   _zz_Array_OUT_227;
  wire       [31:0]   _zz_Array_OUT_228;
  wire       [31:0]   _zz_Array_OUT_229;
  wire       [31:0]   _zz_Array_OUT_230;
  wire       [31:0]   _zz_Array_OUT_231;
  wire       [31:0]   _zz_Array_OUT_232;
  wire       [31:0]   _zz_Array_OUT_233;
  wire       [31:0]   _zz_Array_OUT_234;
  wire       [31:0]   _zz_Array_OUT_235;
  wire       [31:0]   _zz_Array_OUT_236;
  wire       [31:0]   _zz_Array_OUT_237;
  wire       [31:0]   _zz_Array_OUT_238;
  wire       [31:0]   _zz_Array_OUT_239;
  wire       [31:0]   _zz_Array_OUT_240;
  wire       [31:0]   _zz_Array_OUT_241;
  wire       [31:0]   _zz_Array_OUT_242;
  wire       [31:0]   _zz_Array_OUT_243;
  wire       [31:0]   _zz_Array_OUT_244;
  wire       [31:0]   _zz_Array_OUT_245;
  wire       [31:0]   _zz_Array_OUT_246;
  wire       [31:0]   _zz_Array_OUT_247;
  wire       [31:0]   _zz_Array_OUT_248;
  wire       [31:0]   _zz_Array_OUT_249;
  wire       [31:0]   _zz_Array_OUT_250;
  wire       [31:0]   _zz_Array_OUT_251;
  wire       [31:0]   _zz_Array_OUT_252;
  wire       [31:0]   _zz_Array_OUT_253;
  wire       [31:0]   _zz_Array_OUT_254;
  wire       [31:0]   _zz_Array_OUT_255;
  wire       [31:0]   _zz_Array_OUT_256;
  wire       [31:0]   _zz_Array_OUT_257;
  wire       [31:0]   _zz_Array_OUT_258;
  wire       [31:0]   _zz_Array_OUT_259;
  wire       [31:0]   _zz_Array_OUT_260;
  wire       [31:0]   _zz_Array_OUT_261;
  wire       [31:0]   _zz_Array_OUT_262;
  wire       [31:0]   _zz_Array_OUT_263;
  wire       [31:0]   _zz_Array_OUT_264;
  wire       [31:0]   _zz_Array_OUT_265;
  wire       [31:0]   _zz_Array_OUT_266;
  wire       [31:0]   _zz_Array_OUT_267;
  wire       [31:0]   _zz_Array_OUT_268;
  wire       [31:0]   _zz_Array_OUT_269;
  wire       [31:0]   _zz_Array_OUT_270;
  wire       [31:0]   _zz_Array_OUT_271;
  wire       [31:0]   _zz_Array_OUT_272;
  wire       [31:0]   _zz_Array_OUT_273;
  wire       [31:0]   _zz_Array_OUT_274;
  wire       [31:0]   _zz_Array_OUT_275;
  wire       [31:0]   _zz_Array_OUT_276;
  wire       [31:0]   _zz_Array_OUT_277;
  wire       [31:0]   _zz_Array_OUT_278;
  wire       [31:0]   _zz_Array_OUT_279;
  wire       [31:0]   _zz_Array_OUT_280;
  wire       [31:0]   _zz_Array_OUT_281;
  wire       [31:0]   _zz_Array_OUT_282;
  wire       [31:0]   _zz_Array_OUT_283;
  wire       [31:0]   _zz_Array_OUT_284;
  wire       [31:0]   _zz_Array_OUT_285;
  wire       [31:0]   _zz_Array_OUT_286;
  wire       [31:0]   _zz_Array_OUT_287;
  wire       [31:0]   _zz_Array_OUT_288;
  wire       [31:0]   _zz_Array_OUT_289;
  wire       [31:0]   _zz_Array_OUT_290;
  wire       [31:0]   _zz_Array_OUT_291;
  wire       [31:0]   _zz_Array_OUT_292;
  wire       [31:0]   _zz_Array_OUT_293;
  wire       [31:0]   _zz_Array_OUT_294;
  wire       [31:0]   _zz_Array_OUT_295;
  wire       [31:0]   _zz_Array_OUT_296;
  wire       [31:0]   _zz_Array_OUT_297;
  wire       [31:0]   _zz_Array_OUT_298;
  wire       [31:0]   _zz_Array_OUT_299;
  wire       [31:0]   _zz_Array_OUT_300;
  wire       [31:0]   _zz_Array_OUT_301;
  wire       [31:0]   _zz_Array_OUT_302;
  wire       [31:0]   _zz_Array_OUT_303;
  wire       [31:0]   _zz_Array_OUT_304;
  wire       [31:0]   _zz_Array_OUT_305;
  wire       [31:0]   _zz_Array_OUT_306;
  wire       [31:0]   _zz_Array_OUT_307;
  wire       [31:0]   _zz_Array_OUT_308;
  wire       [31:0]   _zz_Array_OUT_309;
  wire       [31:0]   _zz_Array_OUT_310;
  wire       [31:0]   _zz_Array_OUT_311;
  wire       [31:0]   _zz_Array_OUT_312;
  wire       [31:0]   _zz_Array_OUT_313;
  wire       [31:0]   _zz_Array_OUT_314;
  wire       [31:0]   _zz_Array_OUT_315;
  wire       [31:0]   _zz_Array_OUT_316;
  wire       [31:0]   _zz_Array_OUT_317;
  wire       [31:0]   _zz_Array_OUT_318;
  wire       [31:0]   _zz_Array_OUT_319;
  wire       [31:0]   _zz_Array_OUT_320;
  wire       [31:0]   _zz_Array_OUT_321;
  wire       [31:0]   _zz_Array_OUT_322;
  wire       [31:0]   _zz_Array_OUT_323;
  wire       [31:0]   _zz_Array_OUT_324;
  wire       [31:0]   _zz_Array_OUT_325;
  wire       [31:0]   _zz_Array_OUT_326;
  wire       [31:0]   _zz_Array_OUT_327;
  wire       [31:0]   _zz_Array_OUT_328;
  wire       [31:0]   _zz_Array_OUT_329;
  wire       [31:0]   _zz_Array_OUT_330;
  wire       [31:0]   _zz_Array_OUT_331;
  wire       [31:0]   _zz_Array_OUT_332;
  wire       [31:0]   _zz_Array_OUT_333;
  wire       [31:0]   _zz_Array_OUT_334;
  wire       [31:0]   _zz_Array_OUT_335;
  wire       [31:0]   _zz_Array_OUT_336;
  wire       [31:0]   _zz_Array_OUT_337;
  wire       [31:0]   _zz_Array_OUT_338;
  wire       [31:0]   _zz_Array_OUT_339;
  wire       [31:0]   _zz_Array_OUT_340;
  wire       [31:0]   _zz_Array_OUT_341;
  wire       [31:0]   _zz_Array_OUT_342;
  wire       [31:0]   _zz_Array_OUT_343;
  wire       [31:0]   _zz_Array_OUT_344;
  wire       [31:0]   _zz_Array_OUT_345;
  wire       [31:0]   _zz_Array_OUT_346;
  wire       [31:0]   _zz_Array_OUT_347;
  wire       [31:0]   _zz_Array_OUT_348;
  wire       [31:0]   _zz_Array_OUT_349;
  wire       [31:0]   _zz_Array_OUT_350;
  wire       [31:0]   _zz_Array_OUT_351;
  wire       [31:0]   _zz_Array_OUT_352;
  wire       [31:0]   _zz_Array_OUT_353;
  wire       [31:0]   _zz_Array_OUT_354;
  wire       [31:0]   _zz_Array_OUT_355;
  wire       [31:0]   _zz_Array_OUT_356;
  wire       [31:0]   _zz_Array_OUT_357;
  wire       [31:0]   _zz_Array_OUT_358;
  wire       [31:0]   _zz_Array_OUT_359;
  wire       [31:0]   _zz_Array_OUT_360;
  wire       [31:0]   _zz_Array_OUT_361;
  wire       [31:0]   _zz_Array_OUT_362;
  wire       [31:0]   _zz_Array_OUT_363;
  wire       [31:0]   _zz_Array_OUT_364;
  wire       [31:0]   _zz_Array_OUT_365;
  wire       [31:0]   _zz_Array_OUT_366;
  wire       [31:0]   _zz_Array_OUT_367;
  wire       [31:0]   _zz_Array_OUT_368;
  wire       [31:0]   _zz_Array_OUT_369;
  wire       [31:0]   _zz_Array_OUT_370;
  wire       [31:0]   _zz_Array_OUT_371;
  wire       [31:0]   _zz_Array_OUT_372;
  wire       [31:0]   _zz_Array_OUT_373;
  wire       [31:0]   _zz_Array_OUT_374;
  wire       [31:0]   _zz_Array_OUT_375;
  wire       [31:0]   _zz_Array_OUT_376;
  wire       [31:0]   _zz_Array_OUT_377;
  wire       [31:0]   _zz_Array_OUT_378;
  wire       [31:0]   _zz_Array_OUT_379;
  wire       [31:0]   _zz_Array_OUT_380;
  wire       [31:0]   _zz_Array_OUT_381;
  wire       [31:0]   _zz_Array_OUT_382;
  wire       [31:0]   _zz_Array_OUT_383;
  wire       [31:0]   _zz_Array_OUT_384;
  wire       [31:0]   _zz_Array_OUT_385;
  wire       [31:0]   _zz_Array_OUT_386;
  wire       [31:0]   _zz_Array_OUT_387;
  wire       [31:0]   _zz_Array_OUT_388;
  wire       [31:0]   _zz_Array_OUT_389;
  wire       [31:0]   _zz_Array_OUT_390;
  wire       [31:0]   _zz_Array_OUT_391;
  wire       [31:0]   _zz_Array_OUT_392;
  wire       [31:0]   _zz_Array_OUT_393;
  wire       [31:0]   _zz_Array_OUT_394;
  wire       [31:0]   _zz_Array_OUT_395;
  wire       [31:0]   _zz_Array_OUT_396;
  wire       [31:0]   _zz_Array_OUT_397;
  wire       [31:0]   _zz_Array_OUT_398;
  wire       [31:0]   _zz_Array_OUT_399;
  wire       [31:0]   _zz_Array_OUT_400;
  wire       [31:0]   _zz_Array_OUT_401;
  wire       [31:0]   _zz_Array_OUT_402;
  wire       [31:0]   _zz_Array_OUT_403;
  wire       [31:0]   _zz_Array_OUT_404;
  wire       [31:0]   _zz_Array_OUT_405;
  wire       [31:0]   _zz_Array_OUT_406;
  wire       [31:0]   _zz_Array_OUT_407;
  wire       [31:0]   _zz_Array_OUT_408;
  wire       [31:0]   _zz_Array_OUT_409;
  wire       [31:0]   _zz_Array_OUT_410;
  wire       [31:0]   _zz_Array_OUT_411;
  wire       [31:0]   _zz_Array_OUT_412;
  wire       [31:0]   _zz_Array_OUT_413;
  wire       [31:0]   _zz_Array_OUT_414;
  wire       [31:0]   _zz_Array_OUT_415;
  wire       [31:0]   _zz_Array_OUT_416;
  wire       [31:0]   _zz_Array_OUT_417;
  wire       [31:0]   _zz_Array_OUT_418;
  wire       [31:0]   _zz_Array_OUT_419;
  wire       [31:0]   _zz_Array_OUT_420;
  wire       [31:0]   _zz_Array_OUT_421;
  wire       [31:0]   _zz_Array_OUT_422;
  wire       [31:0]   _zz_Array_OUT_423;
  wire       [31:0]   _zz_Array_OUT_424;
  wire       [31:0]   _zz_Array_OUT_425;
  wire       [31:0]   _zz_Array_OUT_426;
  wire       [31:0]   _zz_Array_OUT_427;
  wire       [31:0]   _zz_Array_OUT_428;
  wire       [31:0]   _zz_Array_OUT_429;
  wire       [31:0]   _zz_Array_OUT_430;
  wire       [31:0]   _zz_Array_OUT_431;
  wire       [31:0]   _zz_Array_OUT_432;
  wire       [31:0]   _zz_Array_OUT_433;
  wire       [31:0]   _zz_Array_OUT_434;
  wire       [31:0]   _zz_Array_OUT_435;
  wire       [31:0]   _zz_Array_OUT_436;
  wire       [31:0]   _zz_Array_OUT_437;
  wire       [31:0]   _zz_Array_OUT_438;
  wire       [31:0]   _zz_Array_OUT_439;
  wire       [31:0]   _zz_Array_OUT_440;
  wire       [31:0]   _zz_Array_OUT_441;
  wire       [31:0]   _zz_Array_OUT_442;
  wire       [31:0]   _zz_Array_OUT_443;
  wire       [31:0]   _zz_Array_OUT_444;
  wire       [31:0]   _zz_Array_OUT_445;
  wire       [31:0]   _zz_Array_OUT_446;
  wire       [31:0]   _zz_Array_OUT_447;
  wire       [2047:0] Array_temp_0;
  wire       [2047:0] Array_temp_1;
  wire       [2047:0] Array_temp_2;
  wire       [2047:0] Array_temp_3;
  wire       [2047:0] Array_temp_4;
  wire       [2047:0] Array_temp_5;
  wire       [2047:0] Array_temp_6;
  wire       [2047:0] Array_temp_7;
  reg                 SCLR;
  reg                 last1;
  reg                 last2;
  reg                 CE;
  wire                add_en;
  reg        [14:0]   cnt;
  wire                when_SystolicArray_l45;
  wire                when_SystolicArray_l49;
  wire                when_SystolicArray_l55;
  wire                when_SystolicArray_l63;
  wire                when_SystolicArray_l73;
  wire                when_SystolicArray_l85;
  wire                when_SystolicArray_l99;
  wire                when_SystolicArray_l115;
  wire                when_SystolicArray_l133;
  wire                when_SystolicArray_l149;
  wire                when_SystolicArray_l163;
  wire                when_SystolicArray_l175;
  wire                when_SystolicArray_l185;
  wire                when_SystolicArray_l193;
  wire                when_SystolicArray_l199;

  assign _zz_Array_OUT = (_zz_Array_OUT_1 + Array_temp_7[31 : 0]);
  assign _zz_Array_OUT_1 = (_zz_Array_OUT_2 + Array_temp_6[31 : 0]);
  assign _zz_Array_OUT_2 = (_zz_Array_OUT_3 + Array_temp_5[31 : 0]);
  assign _zz_Array_OUT_3 = (_zz_Array_OUT_4 + Array_temp_4[31 : 0]);
  assign _zz_Array_OUT_4 = (_zz_Array_OUT_5 + Array_temp_3[31 : 0]);
  assign _zz_Array_OUT_5 = (_zz_Array_OUT_6 + Array_temp_2[31 : 0]);
  assign _zz_Array_OUT_6 = (Array_temp_0[31 : 0] + Array_temp_1[31 : 0]);
  assign _zz_Array_OUT_7 = (_zz_Array_OUT_8 + Array_temp_7[63 : 32]);
  assign _zz_Array_OUT_8 = (_zz_Array_OUT_9 + Array_temp_6[63 : 32]);
  assign _zz_Array_OUT_9 = (_zz_Array_OUT_10 + Array_temp_5[63 : 32]);
  assign _zz_Array_OUT_10 = (_zz_Array_OUT_11 + Array_temp_4[63 : 32]);
  assign _zz_Array_OUT_11 = (_zz_Array_OUT_12 + Array_temp_3[63 : 32]);
  assign _zz_Array_OUT_12 = (_zz_Array_OUT_13 + Array_temp_2[63 : 32]);
  assign _zz_Array_OUT_13 = (Array_temp_0[63 : 32] + Array_temp_1[63 : 32]);
  assign _zz_Array_OUT_14 = (_zz_Array_OUT_15 + Array_temp_7[287 : 256]);
  assign _zz_Array_OUT_15 = (_zz_Array_OUT_16 + Array_temp_6[287 : 256]);
  assign _zz_Array_OUT_16 = (_zz_Array_OUT_17 + Array_temp_5[287 : 256]);
  assign _zz_Array_OUT_17 = (_zz_Array_OUT_18 + Array_temp_4[287 : 256]);
  assign _zz_Array_OUT_18 = (_zz_Array_OUT_19 + Array_temp_3[287 : 256]);
  assign _zz_Array_OUT_19 = (_zz_Array_OUT_20 + Array_temp_2[287 : 256]);
  assign _zz_Array_OUT_20 = (Array_temp_0[287 : 256] + Array_temp_1[287 : 256]);
  assign _zz_Array_OUT_21 = (_zz_Array_OUT_22 + Array_temp_7[95 : 64]);
  assign _zz_Array_OUT_22 = (_zz_Array_OUT_23 + Array_temp_6[95 : 64]);
  assign _zz_Array_OUT_23 = (_zz_Array_OUT_24 + Array_temp_5[95 : 64]);
  assign _zz_Array_OUT_24 = (_zz_Array_OUT_25 + Array_temp_4[95 : 64]);
  assign _zz_Array_OUT_25 = (_zz_Array_OUT_26 + Array_temp_3[95 : 64]);
  assign _zz_Array_OUT_26 = (_zz_Array_OUT_27 + Array_temp_2[95 : 64]);
  assign _zz_Array_OUT_27 = (Array_temp_0[95 : 64] + Array_temp_1[95 : 64]);
  assign _zz_Array_OUT_28 = (_zz_Array_OUT_29 + Array_temp_7[543 : 512]);
  assign _zz_Array_OUT_29 = (_zz_Array_OUT_30 + Array_temp_6[543 : 512]);
  assign _zz_Array_OUT_30 = (_zz_Array_OUT_31 + Array_temp_5[543 : 512]);
  assign _zz_Array_OUT_31 = (_zz_Array_OUT_32 + Array_temp_4[543 : 512]);
  assign _zz_Array_OUT_32 = (_zz_Array_OUT_33 + Array_temp_3[543 : 512]);
  assign _zz_Array_OUT_33 = (_zz_Array_OUT_34 + Array_temp_2[543 : 512]);
  assign _zz_Array_OUT_34 = (Array_temp_0[543 : 512] + Array_temp_1[543 : 512]);
  assign _zz_Array_OUT_35 = (_zz_Array_OUT_36 + Array_temp_7[319 : 288]);
  assign _zz_Array_OUT_36 = (_zz_Array_OUT_37 + Array_temp_6[319 : 288]);
  assign _zz_Array_OUT_37 = (_zz_Array_OUT_38 + Array_temp_5[319 : 288]);
  assign _zz_Array_OUT_38 = (_zz_Array_OUT_39 + Array_temp_4[319 : 288]);
  assign _zz_Array_OUT_39 = (_zz_Array_OUT_40 + Array_temp_3[319 : 288]);
  assign _zz_Array_OUT_40 = (_zz_Array_OUT_41 + Array_temp_2[319 : 288]);
  assign _zz_Array_OUT_41 = (Array_temp_0[319 : 288] + Array_temp_1[319 : 288]);
  assign _zz_Array_OUT_42 = (_zz_Array_OUT_43 + Array_temp_7[127 : 96]);
  assign _zz_Array_OUT_43 = (_zz_Array_OUT_44 + Array_temp_6[127 : 96]);
  assign _zz_Array_OUT_44 = (_zz_Array_OUT_45 + Array_temp_5[127 : 96]);
  assign _zz_Array_OUT_45 = (_zz_Array_OUT_46 + Array_temp_4[127 : 96]);
  assign _zz_Array_OUT_46 = (_zz_Array_OUT_47 + Array_temp_3[127 : 96]);
  assign _zz_Array_OUT_47 = (_zz_Array_OUT_48 + Array_temp_2[127 : 96]);
  assign _zz_Array_OUT_48 = (Array_temp_0[127 : 96] + Array_temp_1[127 : 96]);
  assign _zz_Array_OUT_49 = (_zz_Array_OUT_50 + Array_temp_7[799 : 768]);
  assign _zz_Array_OUT_50 = (_zz_Array_OUT_51 + Array_temp_6[799 : 768]);
  assign _zz_Array_OUT_51 = (_zz_Array_OUT_52 + Array_temp_5[799 : 768]);
  assign _zz_Array_OUT_52 = (_zz_Array_OUT_53 + Array_temp_4[799 : 768]);
  assign _zz_Array_OUT_53 = (_zz_Array_OUT_54 + Array_temp_3[799 : 768]);
  assign _zz_Array_OUT_54 = (_zz_Array_OUT_55 + Array_temp_2[799 : 768]);
  assign _zz_Array_OUT_55 = (Array_temp_0[799 : 768] + Array_temp_1[799 : 768]);
  assign _zz_Array_OUT_56 = (_zz_Array_OUT_57 + Array_temp_7[351 : 320]);
  assign _zz_Array_OUT_57 = (_zz_Array_OUT_58 + Array_temp_6[351 : 320]);
  assign _zz_Array_OUT_58 = (_zz_Array_OUT_59 + Array_temp_5[351 : 320]);
  assign _zz_Array_OUT_59 = (_zz_Array_OUT_60 + Array_temp_4[351 : 320]);
  assign _zz_Array_OUT_60 = (_zz_Array_OUT_61 + Array_temp_3[351 : 320]);
  assign _zz_Array_OUT_61 = (_zz_Array_OUT_62 + Array_temp_2[351 : 320]);
  assign _zz_Array_OUT_62 = (Array_temp_0[351 : 320] + Array_temp_1[351 : 320]);
  assign _zz_Array_OUT_63 = (_zz_Array_OUT_64 + Array_temp_7[575 : 544]);
  assign _zz_Array_OUT_64 = (_zz_Array_OUT_65 + Array_temp_6[575 : 544]);
  assign _zz_Array_OUT_65 = (_zz_Array_OUT_66 + Array_temp_5[575 : 544]);
  assign _zz_Array_OUT_66 = (_zz_Array_OUT_67 + Array_temp_4[575 : 544]);
  assign _zz_Array_OUT_67 = (_zz_Array_OUT_68 + Array_temp_3[575 : 544]);
  assign _zz_Array_OUT_68 = (_zz_Array_OUT_69 + Array_temp_2[575 : 544]);
  assign _zz_Array_OUT_69 = (Array_temp_0[575 : 544] + Array_temp_1[575 : 544]);
  assign _zz_Array_OUT_70 = (_zz_Array_OUT_71 + Array_temp_7[159 : 128]);
  assign _zz_Array_OUT_71 = (_zz_Array_OUT_72 + Array_temp_6[159 : 128]);
  assign _zz_Array_OUT_72 = (_zz_Array_OUT_73 + Array_temp_5[159 : 128]);
  assign _zz_Array_OUT_73 = (_zz_Array_OUT_74 + Array_temp_4[159 : 128]);
  assign _zz_Array_OUT_74 = (_zz_Array_OUT_75 + Array_temp_3[159 : 128]);
  assign _zz_Array_OUT_75 = (_zz_Array_OUT_76 + Array_temp_2[159 : 128]);
  assign _zz_Array_OUT_76 = (Array_temp_0[159 : 128] + Array_temp_1[159 : 128]);
  assign _zz_Array_OUT_77 = (_zz_Array_OUT_78 + Array_temp_7[1055 : 1024]);
  assign _zz_Array_OUT_78 = (_zz_Array_OUT_79 + Array_temp_6[1055 : 1024]);
  assign _zz_Array_OUT_79 = (_zz_Array_OUT_80 + Array_temp_5[1055 : 1024]);
  assign _zz_Array_OUT_80 = (_zz_Array_OUT_81 + Array_temp_4[1055 : 1024]);
  assign _zz_Array_OUT_81 = (_zz_Array_OUT_82 + Array_temp_3[1055 : 1024]);
  assign _zz_Array_OUT_82 = (_zz_Array_OUT_83 + Array_temp_2[1055 : 1024]);
  assign _zz_Array_OUT_83 = (Array_temp_0[1055 : 1024] + Array_temp_1[1055 : 1024]);
  assign _zz_Array_OUT_84 = (_zz_Array_OUT_85 + Array_temp_7[383 : 352]);
  assign _zz_Array_OUT_85 = (_zz_Array_OUT_86 + Array_temp_6[383 : 352]);
  assign _zz_Array_OUT_86 = (_zz_Array_OUT_87 + Array_temp_5[383 : 352]);
  assign _zz_Array_OUT_87 = (_zz_Array_OUT_88 + Array_temp_4[383 : 352]);
  assign _zz_Array_OUT_88 = (_zz_Array_OUT_89 + Array_temp_3[383 : 352]);
  assign _zz_Array_OUT_89 = (_zz_Array_OUT_90 + Array_temp_2[383 : 352]);
  assign _zz_Array_OUT_90 = (Array_temp_0[383 : 352] + Array_temp_1[383 : 352]);
  assign _zz_Array_OUT_91 = (_zz_Array_OUT_92 + Array_temp_7[831 : 800]);
  assign _zz_Array_OUT_92 = (_zz_Array_OUT_93 + Array_temp_6[831 : 800]);
  assign _zz_Array_OUT_93 = (_zz_Array_OUT_94 + Array_temp_5[831 : 800]);
  assign _zz_Array_OUT_94 = (_zz_Array_OUT_95 + Array_temp_4[831 : 800]);
  assign _zz_Array_OUT_95 = (_zz_Array_OUT_96 + Array_temp_3[831 : 800]);
  assign _zz_Array_OUT_96 = (_zz_Array_OUT_97 + Array_temp_2[831 : 800]);
  assign _zz_Array_OUT_97 = (Array_temp_0[831 : 800] + Array_temp_1[831 : 800]);
  assign _zz_Array_OUT_98 = (_zz_Array_OUT_99 + Array_temp_7[607 : 576]);
  assign _zz_Array_OUT_99 = (_zz_Array_OUT_100 + Array_temp_6[607 : 576]);
  assign _zz_Array_OUT_100 = (_zz_Array_OUT_101 + Array_temp_5[607 : 576]);
  assign _zz_Array_OUT_101 = (_zz_Array_OUT_102 + Array_temp_4[607 : 576]);
  assign _zz_Array_OUT_102 = (_zz_Array_OUT_103 + Array_temp_3[607 : 576]);
  assign _zz_Array_OUT_103 = (_zz_Array_OUT_104 + Array_temp_2[607 : 576]);
  assign _zz_Array_OUT_104 = (Array_temp_0[607 : 576] + Array_temp_1[607 : 576]);
  assign _zz_Array_OUT_105 = (_zz_Array_OUT_106 + Array_temp_7[191 : 160]);
  assign _zz_Array_OUT_106 = (_zz_Array_OUT_107 + Array_temp_6[191 : 160]);
  assign _zz_Array_OUT_107 = (_zz_Array_OUT_108 + Array_temp_5[191 : 160]);
  assign _zz_Array_OUT_108 = (_zz_Array_OUT_109 + Array_temp_4[191 : 160]);
  assign _zz_Array_OUT_109 = (_zz_Array_OUT_110 + Array_temp_3[191 : 160]);
  assign _zz_Array_OUT_110 = (_zz_Array_OUT_111 + Array_temp_2[191 : 160]);
  assign _zz_Array_OUT_111 = (Array_temp_0[191 : 160] + Array_temp_1[191 : 160]);
  assign _zz_Array_OUT_112 = (_zz_Array_OUT_113 + Array_temp_7[1311 : 1280]);
  assign _zz_Array_OUT_113 = (_zz_Array_OUT_114 + Array_temp_6[1311 : 1280]);
  assign _zz_Array_OUT_114 = (_zz_Array_OUT_115 + Array_temp_5[1311 : 1280]);
  assign _zz_Array_OUT_115 = (_zz_Array_OUT_116 + Array_temp_4[1311 : 1280]);
  assign _zz_Array_OUT_116 = (_zz_Array_OUT_117 + Array_temp_3[1311 : 1280]);
  assign _zz_Array_OUT_117 = (_zz_Array_OUT_118 + Array_temp_2[1311 : 1280]);
  assign _zz_Array_OUT_118 = (Array_temp_0[1311 : 1280] + Array_temp_1[1311 : 1280]);
  assign _zz_Array_OUT_119 = (_zz_Array_OUT_120 + Array_temp_7[415 : 384]);
  assign _zz_Array_OUT_120 = (_zz_Array_OUT_121 + Array_temp_6[415 : 384]);
  assign _zz_Array_OUT_121 = (_zz_Array_OUT_122 + Array_temp_5[415 : 384]);
  assign _zz_Array_OUT_122 = (_zz_Array_OUT_123 + Array_temp_4[415 : 384]);
  assign _zz_Array_OUT_123 = (_zz_Array_OUT_124 + Array_temp_3[415 : 384]);
  assign _zz_Array_OUT_124 = (_zz_Array_OUT_125 + Array_temp_2[415 : 384]);
  assign _zz_Array_OUT_125 = (Array_temp_0[415 : 384] + Array_temp_1[415 : 384]);
  assign _zz_Array_OUT_126 = (_zz_Array_OUT_127 + Array_temp_7[1087 : 1056]);
  assign _zz_Array_OUT_127 = (_zz_Array_OUT_128 + Array_temp_6[1087 : 1056]);
  assign _zz_Array_OUT_128 = (_zz_Array_OUT_129 + Array_temp_5[1087 : 1056]);
  assign _zz_Array_OUT_129 = (_zz_Array_OUT_130 + Array_temp_4[1087 : 1056]);
  assign _zz_Array_OUT_130 = (_zz_Array_OUT_131 + Array_temp_3[1087 : 1056]);
  assign _zz_Array_OUT_131 = (_zz_Array_OUT_132 + Array_temp_2[1087 : 1056]);
  assign _zz_Array_OUT_132 = (Array_temp_0[1087 : 1056] + Array_temp_1[1087 : 1056]);
  assign _zz_Array_OUT_133 = (_zz_Array_OUT_134 + Array_temp_7[639 : 608]);
  assign _zz_Array_OUT_134 = (_zz_Array_OUT_135 + Array_temp_6[639 : 608]);
  assign _zz_Array_OUT_135 = (_zz_Array_OUT_136 + Array_temp_5[639 : 608]);
  assign _zz_Array_OUT_136 = (_zz_Array_OUT_137 + Array_temp_4[639 : 608]);
  assign _zz_Array_OUT_137 = (_zz_Array_OUT_138 + Array_temp_3[639 : 608]);
  assign _zz_Array_OUT_138 = (_zz_Array_OUT_139 + Array_temp_2[639 : 608]);
  assign _zz_Array_OUT_139 = (Array_temp_0[639 : 608] + Array_temp_1[639 : 608]);
  assign _zz_Array_OUT_140 = (_zz_Array_OUT_141 + Array_temp_7[863 : 832]);
  assign _zz_Array_OUT_141 = (_zz_Array_OUT_142 + Array_temp_6[863 : 832]);
  assign _zz_Array_OUT_142 = (_zz_Array_OUT_143 + Array_temp_5[863 : 832]);
  assign _zz_Array_OUT_143 = (_zz_Array_OUT_144 + Array_temp_4[863 : 832]);
  assign _zz_Array_OUT_144 = (_zz_Array_OUT_145 + Array_temp_3[863 : 832]);
  assign _zz_Array_OUT_145 = (_zz_Array_OUT_146 + Array_temp_2[863 : 832]);
  assign _zz_Array_OUT_146 = (Array_temp_0[863 : 832] + Array_temp_1[863 : 832]);
  assign _zz_Array_OUT_147 = (_zz_Array_OUT_148 + Array_temp_7[223 : 192]);
  assign _zz_Array_OUT_148 = (_zz_Array_OUT_149 + Array_temp_6[223 : 192]);
  assign _zz_Array_OUT_149 = (_zz_Array_OUT_150 + Array_temp_5[223 : 192]);
  assign _zz_Array_OUT_150 = (_zz_Array_OUT_151 + Array_temp_4[223 : 192]);
  assign _zz_Array_OUT_151 = (_zz_Array_OUT_152 + Array_temp_3[223 : 192]);
  assign _zz_Array_OUT_152 = (_zz_Array_OUT_153 + Array_temp_2[223 : 192]);
  assign _zz_Array_OUT_153 = (Array_temp_0[223 : 192] + Array_temp_1[223 : 192]);
  assign _zz_Array_OUT_154 = (_zz_Array_OUT_155 + Array_temp_7[1567 : 1536]);
  assign _zz_Array_OUT_155 = (_zz_Array_OUT_156 + Array_temp_6[1567 : 1536]);
  assign _zz_Array_OUT_156 = (_zz_Array_OUT_157 + Array_temp_5[1567 : 1536]);
  assign _zz_Array_OUT_157 = (_zz_Array_OUT_158 + Array_temp_4[1567 : 1536]);
  assign _zz_Array_OUT_158 = (_zz_Array_OUT_159 + Array_temp_3[1567 : 1536]);
  assign _zz_Array_OUT_159 = (_zz_Array_OUT_160 + Array_temp_2[1567 : 1536]);
  assign _zz_Array_OUT_160 = (Array_temp_0[1567 : 1536] + Array_temp_1[1567 : 1536]);
  assign _zz_Array_OUT_161 = (_zz_Array_OUT_162 + Array_temp_7[447 : 416]);
  assign _zz_Array_OUT_162 = (_zz_Array_OUT_163 + Array_temp_6[447 : 416]);
  assign _zz_Array_OUT_163 = (_zz_Array_OUT_164 + Array_temp_5[447 : 416]);
  assign _zz_Array_OUT_164 = (_zz_Array_OUT_165 + Array_temp_4[447 : 416]);
  assign _zz_Array_OUT_165 = (_zz_Array_OUT_166 + Array_temp_3[447 : 416]);
  assign _zz_Array_OUT_166 = (_zz_Array_OUT_167 + Array_temp_2[447 : 416]);
  assign _zz_Array_OUT_167 = (Array_temp_0[447 : 416] + Array_temp_1[447 : 416]);
  assign _zz_Array_OUT_168 = (_zz_Array_OUT_169 + Array_temp_7[1343 : 1312]);
  assign _zz_Array_OUT_169 = (_zz_Array_OUT_170 + Array_temp_6[1343 : 1312]);
  assign _zz_Array_OUT_170 = (_zz_Array_OUT_171 + Array_temp_5[1343 : 1312]);
  assign _zz_Array_OUT_171 = (_zz_Array_OUT_172 + Array_temp_4[1343 : 1312]);
  assign _zz_Array_OUT_172 = (_zz_Array_OUT_173 + Array_temp_3[1343 : 1312]);
  assign _zz_Array_OUT_173 = (_zz_Array_OUT_174 + Array_temp_2[1343 : 1312]);
  assign _zz_Array_OUT_174 = (Array_temp_0[1343 : 1312] + Array_temp_1[1343 : 1312]);
  assign _zz_Array_OUT_175 = (_zz_Array_OUT_176 + Array_temp_7[671 : 640]);
  assign _zz_Array_OUT_176 = (_zz_Array_OUT_177 + Array_temp_6[671 : 640]);
  assign _zz_Array_OUT_177 = (_zz_Array_OUT_178 + Array_temp_5[671 : 640]);
  assign _zz_Array_OUT_178 = (_zz_Array_OUT_179 + Array_temp_4[671 : 640]);
  assign _zz_Array_OUT_179 = (_zz_Array_OUT_180 + Array_temp_3[671 : 640]);
  assign _zz_Array_OUT_180 = (_zz_Array_OUT_181 + Array_temp_2[671 : 640]);
  assign _zz_Array_OUT_181 = (Array_temp_0[671 : 640] + Array_temp_1[671 : 640]);
  assign _zz_Array_OUT_182 = (_zz_Array_OUT_183 + Array_temp_7[1119 : 1088]);
  assign _zz_Array_OUT_183 = (_zz_Array_OUT_184 + Array_temp_6[1119 : 1088]);
  assign _zz_Array_OUT_184 = (_zz_Array_OUT_185 + Array_temp_5[1119 : 1088]);
  assign _zz_Array_OUT_185 = (_zz_Array_OUT_186 + Array_temp_4[1119 : 1088]);
  assign _zz_Array_OUT_186 = (_zz_Array_OUT_187 + Array_temp_3[1119 : 1088]);
  assign _zz_Array_OUT_187 = (_zz_Array_OUT_188 + Array_temp_2[1119 : 1088]);
  assign _zz_Array_OUT_188 = (Array_temp_0[1119 : 1088] + Array_temp_1[1119 : 1088]);
  assign _zz_Array_OUT_189 = (_zz_Array_OUT_190 + Array_temp_7[895 : 864]);
  assign _zz_Array_OUT_190 = (_zz_Array_OUT_191 + Array_temp_6[895 : 864]);
  assign _zz_Array_OUT_191 = (_zz_Array_OUT_192 + Array_temp_5[895 : 864]);
  assign _zz_Array_OUT_192 = (_zz_Array_OUT_193 + Array_temp_4[895 : 864]);
  assign _zz_Array_OUT_193 = (_zz_Array_OUT_194 + Array_temp_3[895 : 864]);
  assign _zz_Array_OUT_194 = (_zz_Array_OUT_195 + Array_temp_2[895 : 864]);
  assign _zz_Array_OUT_195 = (Array_temp_0[895 : 864] + Array_temp_1[895 : 864]);
  assign _zz_Array_OUT_196 = (_zz_Array_OUT_197 + Array_temp_7[255 : 224]);
  assign _zz_Array_OUT_197 = (_zz_Array_OUT_198 + Array_temp_6[255 : 224]);
  assign _zz_Array_OUT_198 = (_zz_Array_OUT_199 + Array_temp_5[255 : 224]);
  assign _zz_Array_OUT_199 = (_zz_Array_OUT_200 + Array_temp_4[255 : 224]);
  assign _zz_Array_OUT_200 = (_zz_Array_OUT_201 + Array_temp_3[255 : 224]);
  assign _zz_Array_OUT_201 = (_zz_Array_OUT_202 + Array_temp_2[255 : 224]);
  assign _zz_Array_OUT_202 = (Array_temp_0[255 : 224] + Array_temp_1[255 : 224]);
  assign _zz_Array_OUT_203 = (_zz_Array_OUT_204 + Array_temp_7[1823 : 1792]);
  assign _zz_Array_OUT_204 = (_zz_Array_OUT_205 + Array_temp_6[1823 : 1792]);
  assign _zz_Array_OUT_205 = (_zz_Array_OUT_206 + Array_temp_5[1823 : 1792]);
  assign _zz_Array_OUT_206 = (_zz_Array_OUT_207 + Array_temp_4[1823 : 1792]);
  assign _zz_Array_OUT_207 = (_zz_Array_OUT_208 + Array_temp_3[1823 : 1792]);
  assign _zz_Array_OUT_208 = (_zz_Array_OUT_209 + Array_temp_2[1823 : 1792]);
  assign _zz_Array_OUT_209 = (Array_temp_0[1823 : 1792] + Array_temp_1[1823 : 1792]);
  assign _zz_Array_OUT_210 = (_zz_Array_OUT_211 + Array_temp_7[479 : 448]);
  assign _zz_Array_OUT_211 = (_zz_Array_OUT_212 + Array_temp_6[479 : 448]);
  assign _zz_Array_OUT_212 = (_zz_Array_OUT_213 + Array_temp_5[479 : 448]);
  assign _zz_Array_OUT_213 = (_zz_Array_OUT_214 + Array_temp_4[479 : 448]);
  assign _zz_Array_OUT_214 = (_zz_Array_OUT_215 + Array_temp_3[479 : 448]);
  assign _zz_Array_OUT_215 = (_zz_Array_OUT_216 + Array_temp_2[479 : 448]);
  assign _zz_Array_OUT_216 = (Array_temp_0[479 : 448] + Array_temp_1[479 : 448]);
  assign _zz_Array_OUT_217 = (_zz_Array_OUT_218 + Array_temp_7[1599 : 1568]);
  assign _zz_Array_OUT_218 = (_zz_Array_OUT_219 + Array_temp_6[1599 : 1568]);
  assign _zz_Array_OUT_219 = (_zz_Array_OUT_220 + Array_temp_5[1599 : 1568]);
  assign _zz_Array_OUT_220 = (_zz_Array_OUT_221 + Array_temp_4[1599 : 1568]);
  assign _zz_Array_OUT_221 = (_zz_Array_OUT_222 + Array_temp_3[1599 : 1568]);
  assign _zz_Array_OUT_222 = (_zz_Array_OUT_223 + Array_temp_2[1599 : 1568]);
  assign _zz_Array_OUT_223 = (Array_temp_0[1599 : 1568] + Array_temp_1[1599 : 1568]);
  assign _zz_Array_OUT_224 = (_zz_Array_OUT_225 + Array_temp_7[703 : 672]);
  assign _zz_Array_OUT_225 = (_zz_Array_OUT_226 + Array_temp_6[703 : 672]);
  assign _zz_Array_OUT_226 = (_zz_Array_OUT_227 + Array_temp_5[703 : 672]);
  assign _zz_Array_OUT_227 = (_zz_Array_OUT_228 + Array_temp_4[703 : 672]);
  assign _zz_Array_OUT_228 = (_zz_Array_OUT_229 + Array_temp_3[703 : 672]);
  assign _zz_Array_OUT_229 = (_zz_Array_OUT_230 + Array_temp_2[703 : 672]);
  assign _zz_Array_OUT_230 = (Array_temp_0[703 : 672] + Array_temp_1[703 : 672]);
  assign _zz_Array_OUT_231 = (_zz_Array_OUT_232 + Array_temp_7[1375 : 1344]);
  assign _zz_Array_OUT_232 = (_zz_Array_OUT_233 + Array_temp_6[1375 : 1344]);
  assign _zz_Array_OUT_233 = (_zz_Array_OUT_234 + Array_temp_5[1375 : 1344]);
  assign _zz_Array_OUT_234 = (_zz_Array_OUT_235 + Array_temp_4[1375 : 1344]);
  assign _zz_Array_OUT_235 = (_zz_Array_OUT_236 + Array_temp_3[1375 : 1344]);
  assign _zz_Array_OUT_236 = (_zz_Array_OUT_237 + Array_temp_2[1375 : 1344]);
  assign _zz_Array_OUT_237 = (Array_temp_0[1375 : 1344] + Array_temp_1[1375 : 1344]);
  assign _zz_Array_OUT_238 = (_zz_Array_OUT_239 + Array_temp_7[927 : 896]);
  assign _zz_Array_OUT_239 = (_zz_Array_OUT_240 + Array_temp_6[927 : 896]);
  assign _zz_Array_OUT_240 = (_zz_Array_OUT_241 + Array_temp_5[927 : 896]);
  assign _zz_Array_OUT_241 = (_zz_Array_OUT_242 + Array_temp_4[927 : 896]);
  assign _zz_Array_OUT_242 = (_zz_Array_OUT_243 + Array_temp_3[927 : 896]);
  assign _zz_Array_OUT_243 = (_zz_Array_OUT_244 + Array_temp_2[927 : 896]);
  assign _zz_Array_OUT_244 = (Array_temp_0[927 : 896] + Array_temp_1[927 : 896]);
  assign _zz_Array_OUT_245 = (_zz_Array_OUT_246 + Array_temp_7[1151 : 1120]);
  assign _zz_Array_OUT_246 = (_zz_Array_OUT_247 + Array_temp_6[1151 : 1120]);
  assign _zz_Array_OUT_247 = (_zz_Array_OUT_248 + Array_temp_5[1151 : 1120]);
  assign _zz_Array_OUT_248 = (_zz_Array_OUT_249 + Array_temp_4[1151 : 1120]);
  assign _zz_Array_OUT_249 = (_zz_Array_OUT_250 + Array_temp_3[1151 : 1120]);
  assign _zz_Array_OUT_250 = (_zz_Array_OUT_251 + Array_temp_2[1151 : 1120]);
  assign _zz_Array_OUT_251 = (Array_temp_0[1151 : 1120] + Array_temp_1[1151 : 1120]);
  assign _zz_Array_OUT_252 = (_zz_Array_OUT_253 + Array_temp_7[511 : 480]);
  assign _zz_Array_OUT_253 = (_zz_Array_OUT_254 + Array_temp_6[511 : 480]);
  assign _zz_Array_OUT_254 = (_zz_Array_OUT_255 + Array_temp_5[511 : 480]);
  assign _zz_Array_OUT_255 = (_zz_Array_OUT_256 + Array_temp_4[511 : 480]);
  assign _zz_Array_OUT_256 = (_zz_Array_OUT_257 + Array_temp_3[511 : 480]);
  assign _zz_Array_OUT_257 = (_zz_Array_OUT_258 + Array_temp_2[511 : 480]);
  assign _zz_Array_OUT_258 = (Array_temp_0[511 : 480] + Array_temp_1[511 : 480]);
  assign _zz_Array_OUT_259 = (_zz_Array_OUT_260 + Array_temp_7[735 : 704]);
  assign _zz_Array_OUT_260 = (_zz_Array_OUT_261 + Array_temp_6[735 : 704]);
  assign _zz_Array_OUT_261 = (_zz_Array_OUT_262 + Array_temp_5[735 : 704]);
  assign _zz_Array_OUT_262 = (_zz_Array_OUT_263 + Array_temp_4[735 : 704]);
  assign _zz_Array_OUT_263 = (_zz_Array_OUT_264 + Array_temp_3[735 : 704]);
  assign _zz_Array_OUT_264 = (_zz_Array_OUT_265 + Array_temp_2[735 : 704]);
  assign _zz_Array_OUT_265 = (Array_temp_0[735 : 704] + Array_temp_1[735 : 704]);
  assign _zz_Array_OUT_266 = (_zz_Array_OUT_267 + Array_temp_7[959 : 928]);
  assign _zz_Array_OUT_267 = (_zz_Array_OUT_268 + Array_temp_6[959 : 928]);
  assign _zz_Array_OUT_268 = (_zz_Array_OUT_269 + Array_temp_5[959 : 928]);
  assign _zz_Array_OUT_269 = (_zz_Array_OUT_270 + Array_temp_4[959 : 928]);
  assign _zz_Array_OUT_270 = (_zz_Array_OUT_271 + Array_temp_3[959 : 928]);
  assign _zz_Array_OUT_271 = (_zz_Array_OUT_272 + Array_temp_2[959 : 928]);
  assign _zz_Array_OUT_272 = (Array_temp_0[959 : 928] + Array_temp_1[959 : 928]);
  assign _zz_Array_OUT_273 = (_zz_Array_OUT_274 + Array_temp_7[1183 : 1152]);
  assign _zz_Array_OUT_274 = (_zz_Array_OUT_275 + Array_temp_6[1183 : 1152]);
  assign _zz_Array_OUT_275 = (_zz_Array_OUT_276 + Array_temp_5[1183 : 1152]);
  assign _zz_Array_OUT_276 = (_zz_Array_OUT_277 + Array_temp_4[1183 : 1152]);
  assign _zz_Array_OUT_277 = (_zz_Array_OUT_278 + Array_temp_3[1183 : 1152]);
  assign _zz_Array_OUT_278 = (_zz_Array_OUT_279 + Array_temp_2[1183 : 1152]);
  assign _zz_Array_OUT_279 = (Array_temp_0[1183 : 1152] + Array_temp_1[1183 : 1152]);
  assign _zz_Array_OUT_280 = (_zz_Array_OUT_281 + Array_temp_7[1407 : 1376]);
  assign _zz_Array_OUT_281 = (_zz_Array_OUT_282 + Array_temp_6[1407 : 1376]);
  assign _zz_Array_OUT_282 = (_zz_Array_OUT_283 + Array_temp_5[1407 : 1376]);
  assign _zz_Array_OUT_283 = (_zz_Array_OUT_284 + Array_temp_4[1407 : 1376]);
  assign _zz_Array_OUT_284 = (_zz_Array_OUT_285 + Array_temp_3[1407 : 1376]);
  assign _zz_Array_OUT_285 = (_zz_Array_OUT_286 + Array_temp_2[1407 : 1376]);
  assign _zz_Array_OUT_286 = (Array_temp_0[1407 : 1376] + Array_temp_1[1407 : 1376]);
  assign _zz_Array_OUT_287 = (_zz_Array_OUT_288 + Array_temp_7[1631 : 1600]);
  assign _zz_Array_OUT_288 = (_zz_Array_OUT_289 + Array_temp_6[1631 : 1600]);
  assign _zz_Array_OUT_289 = (_zz_Array_OUT_290 + Array_temp_5[1631 : 1600]);
  assign _zz_Array_OUT_290 = (_zz_Array_OUT_291 + Array_temp_4[1631 : 1600]);
  assign _zz_Array_OUT_291 = (_zz_Array_OUT_292 + Array_temp_3[1631 : 1600]);
  assign _zz_Array_OUT_292 = (_zz_Array_OUT_293 + Array_temp_2[1631 : 1600]);
  assign _zz_Array_OUT_293 = (Array_temp_0[1631 : 1600] + Array_temp_1[1631 : 1600]);
  assign _zz_Array_OUT_294 = (_zz_Array_OUT_295 + Array_temp_7[1855 : 1824]);
  assign _zz_Array_OUT_295 = (_zz_Array_OUT_296 + Array_temp_6[1855 : 1824]);
  assign _zz_Array_OUT_296 = (_zz_Array_OUT_297 + Array_temp_5[1855 : 1824]);
  assign _zz_Array_OUT_297 = (_zz_Array_OUT_298 + Array_temp_4[1855 : 1824]);
  assign _zz_Array_OUT_298 = (_zz_Array_OUT_299 + Array_temp_3[1855 : 1824]);
  assign _zz_Array_OUT_299 = (_zz_Array_OUT_300 + Array_temp_2[1855 : 1824]);
  assign _zz_Array_OUT_300 = (Array_temp_0[1855 : 1824] + Array_temp_1[1855 : 1824]);
  assign _zz_Array_OUT_301 = (_zz_Array_OUT_302 + Array_temp_7[767 : 736]);
  assign _zz_Array_OUT_302 = (_zz_Array_OUT_303 + Array_temp_6[767 : 736]);
  assign _zz_Array_OUT_303 = (_zz_Array_OUT_304 + Array_temp_5[767 : 736]);
  assign _zz_Array_OUT_304 = (_zz_Array_OUT_305 + Array_temp_4[767 : 736]);
  assign _zz_Array_OUT_305 = (_zz_Array_OUT_306 + Array_temp_3[767 : 736]);
  assign _zz_Array_OUT_306 = (_zz_Array_OUT_307 + Array_temp_2[767 : 736]);
  assign _zz_Array_OUT_307 = (Array_temp_0[767 : 736] + Array_temp_1[767 : 736]);
  assign _zz_Array_OUT_308 = (_zz_Array_OUT_309 + Array_temp_7[991 : 960]);
  assign _zz_Array_OUT_309 = (_zz_Array_OUT_310 + Array_temp_6[991 : 960]);
  assign _zz_Array_OUT_310 = (_zz_Array_OUT_311 + Array_temp_5[991 : 960]);
  assign _zz_Array_OUT_311 = (_zz_Array_OUT_312 + Array_temp_4[991 : 960]);
  assign _zz_Array_OUT_312 = (_zz_Array_OUT_313 + Array_temp_3[991 : 960]);
  assign _zz_Array_OUT_313 = (_zz_Array_OUT_314 + Array_temp_2[991 : 960]);
  assign _zz_Array_OUT_314 = (Array_temp_0[991 : 960] + Array_temp_1[991 : 960]);
  assign _zz_Array_OUT_315 = (_zz_Array_OUT_316 + Array_temp_7[1215 : 1184]);
  assign _zz_Array_OUT_316 = (_zz_Array_OUT_317 + Array_temp_6[1215 : 1184]);
  assign _zz_Array_OUT_317 = (_zz_Array_OUT_318 + Array_temp_5[1215 : 1184]);
  assign _zz_Array_OUT_318 = (_zz_Array_OUT_319 + Array_temp_4[1215 : 1184]);
  assign _zz_Array_OUT_319 = (_zz_Array_OUT_320 + Array_temp_3[1215 : 1184]);
  assign _zz_Array_OUT_320 = (_zz_Array_OUT_321 + Array_temp_2[1215 : 1184]);
  assign _zz_Array_OUT_321 = (Array_temp_0[1215 : 1184] + Array_temp_1[1215 : 1184]);
  assign _zz_Array_OUT_322 = (_zz_Array_OUT_323 + Array_temp_7[1439 : 1408]);
  assign _zz_Array_OUT_323 = (_zz_Array_OUT_324 + Array_temp_6[1439 : 1408]);
  assign _zz_Array_OUT_324 = (_zz_Array_OUT_325 + Array_temp_5[1439 : 1408]);
  assign _zz_Array_OUT_325 = (_zz_Array_OUT_326 + Array_temp_4[1439 : 1408]);
  assign _zz_Array_OUT_326 = (_zz_Array_OUT_327 + Array_temp_3[1439 : 1408]);
  assign _zz_Array_OUT_327 = (_zz_Array_OUT_328 + Array_temp_2[1439 : 1408]);
  assign _zz_Array_OUT_328 = (Array_temp_0[1439 : 1408] + Array_temp_1[1439 : 1408]);
  assign _zz_Array_OUT_329 = (_zz_Array_OUT_330 + Array_temp_7[1663 : 1632]);
  assign _zz_Array_OUT_330 = (_zz_Array_OUT_331 + Array_temp_6[1663 : 1632]);
  assign _zz_Array_OUT_331 = (_zz_Array_OUT_332 + Array_temp_5[1663 : 1632]);
  assign _zz_Array_OUT_332 = (_zz_Array_OUT_333 + Array_temp_4[1663 : 1632]);
  assign _zz_Array_OUT_333 = (_zz_Array_OUT_334 + Array_temp_3[1663 : 1632]);
  assign _zz_Array_OUT_334 = (_zz_Array_OUT_335 + Array_temp_2[1663 : 1632]);
  assign _zz_Array_OUT_335 = (Array_temp_0[1663 : 1632] + Array_temp_1[1663 : 1632]);
  assign _zz_Array_OUT_336 = (_zz_Array_OUT_337 + Array_temp_7[1887 : 1856]);
  assign _zz_Array_OUT_337 = (_zz_Array_OUT_338 + Array_temp_6[1887 : 1856]);
  assign _zz_Array_OUT_338 = (_zz_Array_OUT_339 + Array_temp_5[1887 : 1856]);
  assign _zz_Array_OUT_339 = (_zz_Array_OUT_340 + Array_temp_4[1887 : 1856]);
  assign _zz_Array_OUT_340 = (_zz_Array_OUT_341 + Array_temp_3[1887 : 1856]);
  assign _zz_Array_OUT_341 = (_zz_Array_OUT_342 + Array_temp_2[1887 : 1856]);
  assign _zz_Array_OUT_342 = (Array_temp_0[1887 : 1856] + Array_temp_1[1887 : 1856]);
  assign _zz_Array_OUT_343 = (_zz_Array_OUT_344 + Array_temp_7[1023 : 992]);
  assign _zz_Array_OUT_344 = (_zz_Array_OUT_345 + Array_temp_6[1023 : 992]);
  assign _zz_Array_OUT_345 = (_zz_Array_OUT_346 + Array_temp_5[1023 : 992]);
  assign _zz_Array_OUT_346 = (_zz_Array_OUT_347 + Array_temp_4[1023 : 992]);
  assign _zz_Array_OUT_347 = (_zz_Array_OUT_348 + Array_temp_3[1023 : 992]);
  assign _zz_Array_OUT_348 = (_zz_Array_OUT_349 + Array_temp_2[1023 : 992]);
  assign _zz_Array_OUT_349 = (Array_temp_0[1023 : 992] + Array_temp_1[1023 : 992]);
  assign _zz_Array_OUT_350 = (_zz_Array_OUT_351 + Array_temp_7[1247 : 1216]);
  assign _zz_Array_OUT_351 = (_zz_Array_OUT_352 + Array_temp_6[1247 : 1216]);
  assign _zz_Array_OUT_352 = (_zz_Array_OUT_353 + Array_temp_5[1247 : 1216]);
  assign _zz_Array_OUT_353 = (_zz_Array_OUT_354 + Array_temp_4[1247 : 1216]);
  assign _zz_Array_OUT_354 = (_zz_Array_OUT_355 + Array_temp_3[1247 : 1216]);
  assign _zz_Array_OUT_355 = (_zz_Array_OUT_356 + Array_temp_2[1247 : 1216]);
  assign _zz_Array_OUT_356 = (Array_temp_0[1247 : 1216] + Array_temp_1[1247 : 1216]);
  assign _zz_Array_OUT_357 = (_zz_Array_OUT_358 + Array_temp_7[1471 : 1440]);
  assign _zz_Array_OUT_358 = (_zz_Array_OUT_359 + Array_temp_6[1471 : 1440]);
  assign _zz_Array_OUT_359 = (_zz_Array_OUT_360 + Array_temp_5[1471 : 1440]);
  assign _zz_Array_OUT_360 = (_zz_Array_OUT_361 + Array_temp_4[1471 : 1440]);
  assign _zz_Array_OUT_361 = (_zz_Array_OUT_362 + Array_temp_3[1471 : 1440]);
  assign _zz_Array_OUT_362 = (_zz_Array_OUT_363 + Array_temp_2[1471 : 1440]);
  assign _zz_Array_OUT_363 = (Array_temp_0[1471 : 1440] + Array_temp_1[1471 : 1440]);
  assign _zz_Array_OUT_364 = (_zz_Array_OUT_365 + Array_temp_7[1695 : 1664]);
  assign _zz_Array_OUT_365 = (_zz_Array_OUT_366 + Array_temp_6[1695 : 1664]);
  assign _zz_Array_OUT_366 = (_zz_Array_OUT_367 + Array_temp_5[1695 : 1664]);
  assign _zz_Array_OUT_367 = (_zz_Array_OUT_368 + Array_temp_4[1695 : 1664]);
  assign _zz_Array_OUT_368 = (_zz_Array_OUT_369 + Array_temp_3[1695 : 1664]);
  assign _zz_Array_OUT_369 = (_zz_Array_OUT_370 + Array_temp_2[1695 : 1664]);
  assign _zz_Array_OUT_370 = (Array_temp_0[1695 : 1664] + Array_temp_1[1695 : 1664]);
  assign _zz_Array_OUT_371 = (_zz_Array_OUT_372 + Array_temp_7[1919 : 1888]);
  assign _zz_Array_OUT_372 = (_zz_Array_OUT_373 + Array_temp_6[1919 : 1888]);
  assign _zz_Array_OUT_373 = (_zz_Array_OUT_374 + Array_temp_5[1919 : 1888]);
  assign _zz_Array_OUT_374 = (_zz_Array_OUT_375 + Array_temp_4[1919 : 1888]);
  assign _zz_Array_OUT_375 = (_zz_Array_OUT_376 + Array_temp_3[1919 : 1888]);
  assign _zz_Array_OUT_376 = (_zz_Array_OUT_377 + Array_temp_2[1919 : 1888]);
  assign _zz_Array_OUT_377 = (Array_temp_0[1919 : 1888] + Array_temp_1[1919 : 1888]);
  assign _zz_Array_OUT_378 = (_zz_Array_OUT_379 + Array_temp_7[1279 : 1248]);
  assign _zz_Array_OUT_379 = (_zz_Array_OUT_380 + Array_temp_6[1279 : 1248]);
  assign _zz_Array_OUT_380 = (_zz_Array_OUT_381 + Array_temp_5[1279 : 1248]);
  assign _zz_Array_OUT_381 = (_zz_Array_OUT_382 + Array_temp_4[1279 : 1248]);
  assign _zz_Array_OUT_382 = (_zz_Array_OUT_383 + Array_temp_3[1279 : 1248]);
  assign _zz_Array_OUT_383 = (_zz_Array_OUT_384 + Array_temp_2[1279 : 1248]);
  assign _zz_Array_OUT_384 = (Array_temp_0[1279 : 1248] + Array_temp_1[1279 : 1248]);
  assign _zz_Array_OUT_385 = (_zz_Array_OUT_386 + Array_temp_7[1503 : 1472]);
  assign _zz_Array_OUT_386 = (_zz_Array_OUT_387 + Array_temp_6[1503 : 1472]);
  assign _zz_Array_OUT_387 = (_zz_Array_OUT_388 + Array_temp_5[1503 : 1472]);
  assign _zz_Array_OUT_388 = (_zz_Array_OUT_389 + Array_temp_4[1503 : 1472]);
  assign _zz_Array_OUT_389 = (_zz_Array_OUT_390 + Array_temp_3[1503 : 1472]);
  assign _zz_Array_OUT_390 = (_zz_Array_OUT_391 + Array_temp_2[1503 : 1472]);
  assign _zz_Array_OUT_391 = (Array_temp_0[1503 : 1472] + Array_temp_1[1503 : 1472]);
  assign _zz_Array_OUT_392 = (_zz_Array_OUT_393 + Array_temp_7[1727 : 1696]);
  assign _zz_Array_OUT_393 = (_zz_Array_OUT_394 + Array_temp_6[1727 : 1696]);
  assign _zz_Array_OUT_394 = (_zz_Array_OUT_395 + Array_temp_5[1727 : 1696]);
  assign _zz_Array_OUT_395 = (_zz_Array_OUT_396 + Array_temp_4[1727 : 1696]);
  assign _zz_Array_OUT_396 = (_zz_Array_OUT_397 + Array_temp_3[1727 : 1696]);
  assign _zz_Array_OUT_397 = (_zz_Array_OUT_398 + Array_temp_2[1727 : 1696]);
  assign _zz_Array_OUT_398 = (Array_temp_0[1727 : 1696] + Array_temp_1[1727 : 1696]);
  assign _zz_Array_OUT_399 = (_zz_Array_OUT_400 + Array_temp_7[1951 : 1920]);
  assign _zz_Array_OUT_400 = (_zz_Array_OUT_401 + Array_temp_6[1951 : 1920]);
  assign _zz_Array_OUT_401 = (_zz_Array_OUT_402 + Array_temp_5[1951 : 1920]);
  assign _zz_Array_OUT_402 = (_zz_Array_OUT_403 + Array_temp_4[1951 : 1920]);
  assign _zz_Array_OUT_403 = (_zz_Array_OUT_404 + Array_temp_3[1951 : 1920]);
  assign _zz_Array_OUT_404 = (_zz_Array_OUT_405 + Array_temp_2[1951 : 1920]);
  assign _zz_Array_OUT_405 = (Array_temp_0[1951 : 1920] + Array_temp_1[1951 : 1920]);
  assign _zz_Array_OUT_406 = (_zz_Array_OUT_407 + Array_temp_7[1535 : 1504]);
  assign _zz_Array_OUT_407 = (_zz_Array_OUT_408 + Array_temp_6[1535 : 1504]);
  assign _zz_Array_OUT_408 = (_zz_Array_OUT_409 + Array_temp_5[1535 : 1504]);
  assign _zz_Array_OUT_409 = (_zz_Array_OUT_410 + Array_temp_4[1535 : 1504]);
  assign _zz_Array_OUT_410 = (_zz_Array_OUT_411 + Array_temp_3[1535 : 1504]);
  assign _zz_Array_OUT_411 = (_zz_Array_OUT_412 + Array_temp_2[1535 : 1504]);
  assign _zz_Array_OUT_412 = (Array_temp_0[1535 : 1504] + Array_temp_1[1535 : 1504]);
  assign _zz_Array_OUT_413 = (_zz_Array_OUT_414 + Array_temp_7[1759 : 1728]);
  assign _zz_Array_OUT_414 = (_zz_Array_OUT_415 + Array_temp_6[1759 : 1728]);
  assign _zz_Array_OUT_415 = (_zz_Array_OUT_416 + Array_temp_5[1759 : 1728]);
  assign _zz_Array_OUT_416 = (_zz_Array_OUT_417 + Array_temp_4[1759 : 1728]);
  assign _zz_Array_OUT_417 = (_zz_Array_OUT_418 + Array_temp_3[1759 : 1728]);
  assign _zz_Array_OUT_418 = (_zz_Array_OUT_419 + Array_temp_2[1759 : 1728]);
  assign _zz_Array_OUT_419 = (Array_temp_0[1759 : 1728] + Array_temp_1[1759 : 1728]);
  assign _zz_Array_OUT_420 = (_zz_Array_OUT_421 + Array_temp_7[1983 : 1952]);
  assign _zz_Array_OUT_421 = (_zz_Array_OUT_422 + Array_temp_6[1983 : 1952]);
  assign _zz_Array_OUT_422 = (_zz_Array_OUT_423 + Array_temp_5[1983 : 1952]);
  assign _zz_Array_OUT_423 = (_zz_Array_OUT_424 + Array_temp_4[1983 : 1952]);
  assign _zz_Array_OUT_424 = (_zz_Array_OUT_425 + Array_temp_3[1983 : 1952]);
  assign _zz_Array_OUT_425 = (_zz_Array_OUT_426 + Array_temp_2[1983 : 1952]);
  assign _zz_Array_OUT_426 = (Array_temp_0[1983 : 1952] + Array_temp_1[1983 : 1952]);
  assign _zz_Array_OUT_427 = (_zz_Array_OUT_428 + Array_temp_7[1791 : 1760]);
  assign _zz_Array_OUT_428 = (_zz_Array_OUT_429 + Array_temp_6[1791 : 1760]);
  assign _zz_Array_OUT_429 = (_zz_Array_OUT_430 + Array_temp_5[1791 : 1760]);
  assign _zz_Array_OUT_430 = (_zz_Array_OUT_431 + Array_temp_4[1791 : 1760]);
  assign _zz_Array_OUT_431 = (_zz_Array_OUT_432 + Array_temp_3[1791 : 1760]);
  assign _zz_Array_OUT_432 = (_zz_Array_OUT_433 + Array_temp_2[1791 : 1760]);
  assign _zz_Array_OUT_433 = (Array_temp_0[1791 : 1760] + Array_temp_1[1791 : 1760]);
  assign _zz_Array_OUT_434 = (_zz_Array_OUT_435 + Array_temp_7[2015 : 1984]);
  assign _zz_Array_OUT_435 = (_zz_Array_OUT_436 + Array_temp_6[2015 : 1984]);
  assign _zz_Array_OUT_436 = (_zz_Array_OUT_437 + Array_temp_5[2015 : 1984]);
  assign _zz_Array_OUT_437 = (_zz_Array_OUT_438 + Array_temp_4[2015 : 1984]);
  assign _zz_Array_OUT_438 = (_zz_Array_OUT_439 + Array_temp_3[2015 : 1984]);
  assign _zz_Array_OUT_439 = (_zz_Array_OUT_440 + Array_temp_2[2015 : 1984]);
  assign _zz_Array_OUT_440 = (Array_temp_0[2015 : 1984] + Array_temp_1[2015 : 1984]);
  assign _zz_Array_OUT_441 = (_zz_Array_OUT_442 + Array_temp_7[2047 : 2016]);
  assign _zz_Array_OUT_442 = (_zz_Array_OUT_443 + Array_temp_6[2047 : 2016]);
  assign _zz_Array_OUT_443 = (_zz_Array_OUT_444 + Array_temp_5[2047 : 2016]);
  assign _zz_Array_OUT_444 = (_zz_Array_OUT_445 + Array_temp_4[2047 : 2016]);
  assign _zz_Array_OUT_445 = (_zz_Array_OUT_446 + Array_temp_3[2047 : 2016]);
  assign _zz_Array_OUT_446 = (_zz_Array_OUT_447 + Array_temp_2[2047 : 2016]);
  assign _zz_Array_OUT_447 = (Array_temp_0[2047 : 2016] + Array_temp_1[2047 : 2016]);
  Tile tile_8 (
    .CE       (CE                     ), //i
    .SCLR     (SCLR                   ), //i
    .A        (tile_8_A[63:0]         ), //i
    .B        (tile_8_B[63:0]         ), //i
    .Tile_OUT (tile_8_Tile_OUT[2047:0]), //o
    .clk      (clk                    ), //i
    .reset    (reset                  )  //i
  );
  Tile tile_9 (
    .CE       (CE                     ), //i
    .SCLR     (SCLR                   ), //i
    .A        (tile_9_A[63:0]         ), //i
    .B        (tile_9_B[63:0]         ), //i
    .Tile_OUT (tile_9_Tile_OUT[2047:0]), //o
    .clk      (clk                    ), //i
    .reset    (reset                  )  //i
  );
  Tile tile_10 (
    .CE       (CE                      ), //i
    .SCLR     (SCLR                    ), //i
    .A        (tile_10_A[63:0]         ), //i
    .B        (tile_10_B[63:0]         ), //i
    .Tile_OUT (tile_10_Tile_OUT[2047:0]), //o
    .clk      (clk                     ), //i
    .reset    (reset                   )  //i
  );
  Tile tile_11 (
    .CE       (CE                      ), //i
    .SCLR     (SCLR                    ), //i
    .A        (tile_11_A[63:0]         ), //i
    .B        (tile_11_B[63:0]         ), //i
    .Tile_OUT (tile_11_Tile_OUT[2047:0]), //o
    .clk      (clk                     ), //i
    .reset    (reset                   )  //i
  );
  Tile tile_12 (
    .CE       (CE                      ), //i
    .SCLR     (SCLR                    ), //i
    .A        (tile_12_A[63:0]         ), //i
    .B        (tile_12_B[63:0]         ), //i
    .Tile_OUT (tile_12_Tile_OUT[2047:0]), //o
    .clk      (clk                     ), //i
    .reset    (reset                   )  //i
  );
  Tile tile_13 (
    .CE       (CE                      ), //i
    .SCLR     (SCLR                    ), //i
    .A        (tile_13_A[63:0]         ), //i
    .B        (tile_13_B[63:0]         ), //i
    .Tile_OUT (tile_13_Tile_OUT[2047:0]), //o
    .clk      (clk                     ), //i
    .reset    (reset                   )  //i
  );
  Tile tile_14 (
    .CE       (CE                      ), //i
    .SCLR     (SCLR                    ), //i
    .A        (tile_14_A[63:0]         ), //i
    .B        (tile_14_B[63:0]         ), //i
    .Tile_OUT (tile_14_Tile_OUT[2047:0]), //o
    .clk      (clk                     ), //i
    .reset    (reset                   )  //i
  );
  Tile tile_15 (
    .CE       (CE                      ), //i
    .SCLR     (SCLR                    ), //i
    .A        (tile_15_A[63:0]         ), //i
    .B        (tile_15_B[63:0]         ), //i
    .Tile_OUT (tile_15_Tile_OUT[2047:0]), //o
    .clk      (clk                     ), //i
    .reset    (reset                   )  //i
  );
  assign add_en = 1'b0;
  assign tile_8_A = A_Array[63 : 0];
  assign tile_8_B = B_Array[63 : 0];
  assign Array_temp_0 = tile_8_Tile_OUT;
  assign tile_9_A = A_Array[127 : 64];
  assign tile_9_B = B_Array[127 : 64];
  assign Array_temp_1 = tile_9_Tile_OUT;
  assign tile_10_A = A_Array[191 : 128];
  assign tile_10_B = B_Array[191 : 128];
  assign Array_temp_2 = tile_10_Tile_OUT;
  assign tile_11_A = A_Array[255 : 192];
  assign tile_11_B = B_Array[255 : 192];
  assign Array_temp_3 = tile_11_Tile_OUT;
  assign tile_12_A = A_Array[319 : 256];
  assign tile_12_B = B_Array[319 : 256];
  assign Array_temp_4 = tile_12_Tile_OUT;
  assign tile_13_A = A_Array[383 : 320];
  assign tile_13_B = B_Array[383 : 320];
  assign Array_temp_5 = tile_13_Tile_OUT;
  assign tile_14_A = A_Array[447 : 384];
  assign tile_14_B = B_Array[447 : 384];
  assign Array_temp_6 = tile_14_Tile_OUT;
  assign tile_15_A = A_Array[511 : 448];
  assign tile_15_B = B_Array[511 : 448];
  assign Array_temp_7 = tile_15_Tile_OUT;
  assign when_SystolicArray_l45 = cnt[0];
  always @(*) begin
    if(when_SystolicArray_l45) begin
      Array_OUT = 2048'h0;
      Array_OUT[31 : 0] = _zz_Array_OUT;
    end else begin
      if(when_SystolicArray_l49) begin
        Array_OUT = 2048'h0;
        Array_OUT[63 : 32] = _zz_Array_OUT_7;
        Array_OUT[287 : 256] = _zz_Array_OUT_14;
      end else begin
        if(when_SystolicArray_l55) begin
          Array_OUT = 2048'h0;
          Array_OUT[95 : 64] = _zz_Array_OUT_21;
          Array_OUT[543 : 512] = _zz_Array_OUT_28;
          Array_OUT[319 : 288] = _zz_Array_OUT_35;
        end else begin
          if(when_SystolicArray_l63) begin
            Array_OUT = 2048'h0;
            Array_OUT[127 : 96] = _zz_Array_OUT_42;
            Array_OUT[799 : 768] = _zz_Array_OUT_49;
            Array_OUT[351 : 320] = _zz_Array_OUT_56;
            Array_OUT[575 : 544] = _zz_Array_OUT_63;
          end else begin
            if(when_SystolicArray_l73) begin
              Array_OUT = 2048'h0;
              Array_OUT[159 : 128] = _zz_Array_OUT_70;
              Array_OUT[1055 : 1024] = _zz_Array_OUT_77;
              Array_OUT[383 : 352] = _zz_Array_OUT_84;
              Array_OUT[831 : 800] = _zz_Array_OUT_91;
              Array_OUT[607 : 576] = _zz_Array_OUT_98;
            end else begin
              if(when_SystolicArray_l85) begin
                Array_OUT = 2048'h0;
                Array_OUT[191 : 160] = _zz_Array_OUT_105;
                Array_OUT[1311 : 1280] = _zz_Array_OUT_112;
                Array_OUT[415 : 384] = _zz_Array_OUT_119;
                Array_OUT[1087 : 1056] = _zz_Array_OUT_126;
                Array_OUT[639 : 608] = _zz_Array_OUT_133;
                Array_OUT[863 : 832] = _zz_Array_OUT_140;
              end else begin
                if(when_SystolicArray_l99) begin
                  Array_OUT = 2048'h0;
                  Array_OUT[223 : 192] = _zz_Array_OUT_147;
                  Array_OUT[1567 : 1536] = _zz_Array_OUT_154;
                  Array_OUT[447 : 416] = _zz_Array_OUT_161;
                  Array_OUT[1343 : 1312] = _zz_Array_OUT_168;
                  Array_OUT[671 : 640] = _zz_Array_OUT_175;
                  Array_OUT[1119 : 1088] = _zz_Array_OUT_182;
                  Array_OUT[895 : 864] = _zz_Array_OUT_189;
                end else begin
                  if(when_SystolicArray_l115) begin
                    Array_OUT = 2048'h0;
                    Array_OUT[255 : 224] = _zz_Array_OUT_196;
                    Array_OUT[1823 : 1792] = _zz_Array_OUT_203;
                    Array_OUT[479 : 448] = _zz_Array_OUT_210;
                    Array_OUT[1599 : 1568] = _zz_Array_OUT_217;
                    Array_OUT[703 : 672] = _zz_Array_OUT_224;
                    Array_OUT[1375 : 1344] = _zz_Array_OUT_231;
                    Array_OUT[927 : 896] = _zz_Array_OUT_238;
                    Array_OUT[1151 : 1120] = _zz_Array_OUT_245;
                  end else begin
                    if(when_SystolicArray_l133) begin
                      Array_OUT = 2048'h0;
                      Array_OUT[511 : 480] = _zz_Array_OUT_252;
                      Array_OUT[735 : 704] = _zz_Array_OUT_259;
                      Array_OUT[959 : 928] = _zz_Array_OUT_266;
                      Array_OUT[1183 : 1152] = _zz_Array_OUT_273;
                      Array_OUT[1407 : 1376] = _zz_Array_OUT_280;
                      Array_OUT[1631 : 1600] = _zz_Array_OUT_287;
                      Array_OUT[1855 : 1824] = _zz_Array_OUT_294;
                    end else begin
                      if(when_SystolicArray_l149) begin
                        Array_OUT = 2048'h0;
                        Array_OUT[767 : 736] = _zz_Array_OUT_301;
                        Array_OUT[991 : 960] = _zz_Array_OUT_308;
                        Array_OUT[1215 : 1184] = _zz_Array_OUT_315;
                        Array_OUT[1439 : 1408] = _zz_Array_OUT_322;
                        Array_OUT[1663 : 1632] = _zz_Array_OUT_329;
                        Array_OUT[1887 : 1856] = _zz_Array_OUT_336;
                      end else begin
                        if(when_SystolicArray_l163) begin
                          Array_OUT = 2048'h0;
                          Array_OUT[1023 : 992] = _zz_Array_OUT_343;
                          Array_OUT[1247 : 1216] = _zz_Array_OUT_350;
                          Array_OUT[1471 : 1440] = _zz_Array_OUT_357;
                          Array_OUT[1695 : 1664] = _zz_Array_OUT_364;
                          Array_OUT[1919 : 1888] = _zz_Array_OUT_371;
                        end else begin
                          if(when_SystolicArray_l175) begin
                            Array_OUT = 2048'h0;
                            Array_OUT[1279 : 1248] = _zz_Array_OUT_378;
                            Array_OUT[1503 : 1472] = _zz_Array_OUT_385;
                            Array_OUT[1727 : 1696] = _zz_Array_OUT_392;
                            Array_OUT[1951 : 1920] = _zz_Array_OUT_399;
                          end else begin
                            if(when_SystolicArray_l185) begin
                              Array_OUT = 2048'h0;
                              Array_OUT[1535 : 1504] = _zz_Array_OUT_406;
                              Array_OUT[1759 : 1728] = _zz_Array_OUT_413;
                              Array_OUT[1983 : 1952] = _zz_Array_OUT_420;
                            end else begin
                              if(when_SystolicArray_l193) begin
                                Array_OUT = 2048'h0;
                                Array_OUT[1791 : 1760] = _zz_Array_OUT_427;
                                Array_OUT[2015 : 1984] = _zz_Array_OUT_434;
                              end else begin
                                if(when_SystolicArray_l199) begin
                                  Array_OUT = 2048'h0;
                                  Array_OUT[2047 : 2016] = _zz_Array_OUT_441;
                                end else begin
                                  Array_OUT = 2048'h0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end

  assign when_SystolicArray_l49 = cnt[1];
  assign when_SystolicArray_l55 = cnt[2];
  assign when_SystolicArray_l63 = cnt[3];
  assign when_SystolicArray_l73 = cnt[4];
  assign when_SystolicArray_l85 = cnt[5];
  assign when_SystolicArray_l99 = cnt[6];
  assign when_SystolicArray_l115 = cnt[7];
  assign when_SystolicArray_l133 = cnt[8];
  assign when_SystolicArray_l149 = cnt[9];
  assign when_SystolicArray_l163 = cnt[10];
  assign when_SystolicArray_l175 = cnt[11];
  assign when_SystolicArray_l185 = cnt[12];
  assign when_SystolicArray_l193 = cnt[13];
  assign when_SystolicArray_l199 = cnt[14];
  always @(posedge clk) begin
    if(reset) begin
      SCLR <= 1'b0;
      last1 <= 1'b0;
      last2 <= 1'b0;
      CE <= 1'b0;
      cnt <= 15'h0;
    end else begin
      CE <= start;
      last1 <= last;
      last2 <= last1;
      SCLR <= last2;
      cnt[0] <= last2;
      cnt[1] <= cnt[0];
      cnt[2] <= cnt[1];
      cnt[3] <= cnt[2];
      cnt[4] <= cnt[3];
      cnt[5] <= cnt[4];
      cnt[6] <= cnt[5];
      cnt[7] <= cnt[6];
      cnt[8] <= cnt[7];
      cnt[9] <= cnt[8];
      cnt[10] <= cnt[9];
      cnt[11] <= cnt[10];
      cnt[12] <= cnt[11];
      cnt[13] <= cnt[12];
      cnt[14] <= cnt[13];
    end
  end


endmodule

//Tile replaced by Tile

//Tile replaced by Tile

//Tile replaced by Tile

//Tile replaced by Tile

//Tile replaced by Tile

//Tile replaced by Tile

//Tile replaced by Tile

module Tile (
  input               CE,
  input               SCLR,
  input      [63:0]   A,
  input      [63:0]   B,
  output reg [2047:0] Tile_OUT,
  input               clk,
  input               reset
);

  wire       [7:0]    pe_00_a;
  wire       [7:0]    pe_00_b;
  wire                pE_1_CE;
  wire                pE_1_SCLR;
  wire       [7:0]    pE_1_b;
  wire                pE_2_CE;
  wire                pE_2_SCLR;
  wire       [7:0]    pE_2_b;
  wire                pE_3_CE;
  wire                pE_3_SCLR;
  wire       [7:0]    pE_3_b;
  wire                pE_4_CE;
  wire                pE_4_SCLR;
  wire       [7:0]    pE_4_b;
  wire                pE_5_CE;
  wire                pE_5_SCLR;
  wire       [7:0]    pE_5_b;
  wire                pE_6_CE;
  wire                pE_6_SCLR;
  wire       [7:0]    pE_6_b;
  wire                pE_7_CE;
  wire                pE_7_SCLR;
  wire       [7:0]    pE_7_b;
  wire                pE_8_CE;
  wire                pE_8_SCLR;
  wire       [7:0]    pE_8_a;
  wire                pE_9_CE;
  wire                pE_9_SCLR;
  wire       [7:0]    pE_9_a;
  wire                pE_10_CE;
  wire                pE_10_SCLR;
  wire       [7:0]    pE_10_a;
  wire                pE_11_CE;
  wire                pE_11_SCLR;
  wire       [7:0]    pE_11_a;
  wire                pE_12_CE;
  wire                pE_12_SCLR;
  wire       [7:0]    pE_12_a;
  wire                pE_13_CE;
  wire                pE_13_SCLR;
  wire       [7:0]    pE_13_a;
  wire                pE_14_CE;
  wire                pE_14_SCLR;
  wire       [7:0]    pE_14_a;
  wire                pE_15_CE;
  wire                pE_15_SCLR;
  wire                pE_16_CE;
  wire                pE_16_SCLR;
  wire                pE_17_CE;
  wire                pE_17_SCLR;
  wire                pE_18_CE;
  wire                pE_18_SCLR;
  wire                pE_19_CE;
  wire                pE_19_SCLR;
  wire                pE_20_CE;
  wire                pE_20_SCLR;
  wire                pE_21_CE;
  wire                pE_21_SCLR;
  wire                pE_22_CE;
  wire                pE_22_SCLR;
  wire                pE_23_CE;
  wire                pE_23_SCLR;
  wire                pE_24_CE;
  wire                pE_24_SCLR;
  wire                pE_25_CE;
  wire                pE_25_SCLR;
  wire                pE_26_CE;
  wire                pE_26_SCLR;
  wire                pE_27_CE;
  wire                pE_27_SCLR;
  wire                pE_28_CE;
  wire                pE_28_SCLR;
  wire                pE_29_CE;
  wire                pE_29_SCLR;
  wire                pE_30_CE;
  wire                pE_30_SCLR;
  wire                pE_31_CE;
  wire                pE_31_SCLR;
  wire                pE_32_CE;
  wire                pE_32_SCLR;
  wire                pE_33_CE;
  wire                pE_33_SCLR;
  wire                pE_34_CE;
  wire                pE_34_SCLR;
  wire                pE_35_CE;
  wire                pE_35_SCLR;
  wire                pE_36_CE;
  wire                pE_36_SCLR;
  wire                pE_37_CE;
  wire                pE_37_SCLR;
  wire                pE_38_CE;
  wire                pE_38_SCLR;
  wire                pE_39_CE;
  wire                pE_39_SCLR;
  wire                pE_40_CE;
  wire                pE_40_SCLR;
  wire                pE_41_CE;
  wire                pE_41_SCLR;
  wire                pE_42_CE;
  wire                pE_42_SCLR;
  wire                pE_43_CE;
  wire                pE_43_SCLR;
  wire                pE_44_CE;
  wire                pE_44_SCLR;
  wire                pE_45_CE;
  wire                pE_45_SCLR;
  wire                pE_46_CE;
  wire                pE_46_SCLR;
  wire                pE_47_CE;
  wire                pE_47_SCLR;
  wire                pE_48_CE;
  wire                pE_48_SCLR;
  wire                pE_49_CE;
  wire                pE_49_SCLR;
  wire                pE_50_CE;
  wire                pE_50_SCLR;
  wire                pE_51_CE;
  wire                pE_51_SCLR;
  wire                pE_52_CE;
  wire                pE_52_SCLR;
  wire                pE_53_CE;
  wire                pE_53_SCLR;
  wire                pE_54_CE;
  wire                pE_54_SCLR;
  wire                pE_55_CE;
  wire                pE_55_SCLR;
  wire                pE_56_CE;
  wire                pE_56_SCLR;
  wire                pE_57_CE;
  wire                pE_57_SCLR;
  wire                pE_58_CE;
  wire                pE_58_SCLR;
  wire                pE_59_CE;
  wire                pE_59_SCLR;
  wire                pE_60_CE;
  wire                pE_60_SCLR;
  wire                pE_61_CE;
  wire                pE_61_SCLR;
  wire                pE_62_CE;
  wire                pE_62_SCLR;
  wire                pE_63_CE;
  wire                pE_63_SCLR;
  wire       [31:0]   pe_00_pe_out;
  wire       [7:0]    pe_00_acout;
  wire       [7:0]    pe_00_bcout;
  wire       [31:0]   pE_1_pe_out;
  wire       [7:0]    pE_1_acout;
  wire       [7:0]    pE_1_bcout;
  wire       [31:0]   pE_2_pe_out;
  wire       [7:0]    pE_2_acout;
  wire       [7:0]    pE_2_bcout;
  wire       [31:0]   pE_3_pe_out;
  wire       [7:0]    pE_3_acout;
  wire       [7:0]    pE_3_bcout;
  wire       [31:0]   pE_4_pe_out;
  wire       [7:0]    pE_4_acout;
  wire       [7:0]    pE_4_bcout;
  wire       [31:0]   pE_5_pe_out;
  wire       [7:0]    pE_5_acout;
  wire       [7:0]    pE_5_bcout;
  wire       [31:0]   pE_6_pe_out;
  wire       [7:0]    pE_6_acout;
  wire       [7:0]    pE_6_bcout;
  wire       [31:0]   pE_7_pe_out;
  wire       [7:0]    pE_7_acout;
  wire       [7:0]    pE_7_bcout;
  wire       [31:0]   pE_8_pe_out;
  wire       [7:0]    pE_8_acout;
  wire       [7:0]    pE_8_bcout;
  wire       [31:0]   pE_9_pe_out;
  wire       [7:0]    pE_9_acout;
  wire       [7:0]    pE_9_bcout;
  wire       [31:0]   pE_10_pe_out;
  wire       [7:0]    pE_10_acout;
  wire       [7:0]    pE_10_bcout;
  wire       [31:0]   pE_11_pe_out;
  wire       [7:0]    pE_11_acout;
  wire       [7:0]    pE_11_bcout;
  wire       [31:0]   pE_12_pe_out;
  wire       [7:0]    pE_12_acout;
  wire       [7:0]    pE_12_bcout;
  wire       [31:0]   pE_13_pe_out;
  wire       [7:0]    pE_13_acout;
  wire       [7:0]    pE_13_bcout;
  wire       [31:0]   pE_14_pe_out;
  wire       [7:0]    pE_14_acout;
  wire       [7:0]    pE_14_bcout;
  wire       [31:0]   pE_15_pe_out;
  wire       [7:0]    pE_15_acout;
  wire       [7:0]    pE_15_bcout;
  wire       [31:0]   pE_16_pe_out;
  wire       [7:0]    pE_16_acout;
  wire       [7:0]    pE_16_bcout;
  wire       [31:0]   pE_17_pe_out;
  wire       [7:0]    pE_17_acout;
  wire       [7:0]    pE_17_bcout;
  wire       [31:0]   pE_18_pe_out;
  wire       [7:0]    pE_18_acout;
  wire       [7:0]    pE_18_bcout;
  wire       [31:0]   pE_19_pe_out;
  wire       [7:0]    pE_19_acout;
  wire       [7:0]    pE_19_bcout;
  wire       [31:0]   pE_20_pe_out;
  wire       [7:0]    pE_20_acout;
  wire       [7:0]    pE_20_bcout;
  wire       [31:0]   pE_21_pe_out;
  wire       [7:0]    pE_21_acout;
  wire       [7:0]    pE_21_bcout;
  wire       [31:0]   pE_22_pe_out;
  wire       [7:0]    pE_22_acout;
  wire       [7:0]    pE_22_bcout;
  wire       [31:0]   pE_23_pe_out;
  wire       [7:0]    pE_23_acout;
  wire       [7:0]    pE_23_bcout;
  wire       [31:0]   pE_24_pe_out;
  wire       [7:0]    pE_24_acout;
  wire       [7:0]    pE_24_bcout;
  wire       [31:0]   pE_25_pe_out;
  wire       [7:0]    pE_25_acout;
  wire       [7:0]    pE_25_bcout;
  wire       [31:0]   pE_26_pe_out;
  wire       [7:0]    pE_26_acout;
  wire       [7:0]    pE_26_bcout;
  wire       [31:0]   pE_27_pe_out;
  wire       [7:0]    pE_27_acout;
  wire       [7:0]    pE_27_bcout;
  wire       [31:0]   pE_28_pe_out;
  wire       [7:0]    pE_28_acout;
  wire       [7:0]    pE_28_bcout;
  wire       [31:0]   pE_29_pe_out;
  wire       [7:0]    pE_29_acout;
  wire       [7:0]    pE_29_bcout;
  wire       [31:0]   pE_30_pe_out;
  wire       [7:0]    pE_30_acout;
  wire       [7:0]    pE_30_bcout;
  wire       [31:0]   pE_31_pe_out;
  wire       [7:0]    pE_31_acout;
  wire       [7:0]    pE_31_bcout;
  wire       [31:0]   pE_32_pe_out;
  wire       [7:0]    pE_32_acout;
  wire       [7:0]    pE_32_bcout;
  wire       [31:0]   pE_33_pe_out;
  wire       [7:0]    pE_33_acout;
  wire       [7:0]    pE_33_bcout;
  wire       [31:0]   pE_34_pe_out;
  wire       [7:0]    pE_34_acout;
  wire       [7:0]    pE_34_bcout;
  wire       [31:0]   pE_35_pe_out;
  wire       [7:0]    pE_35_acout;
  wire       [7:0]    pE_35_bcout;
  wire       [31:0]   pE_36_pe_out;
  wire       [7:0]    pE_36_acout;
  wire       [7:0]    pE_36_bcout;
  wire       [31:0]   pE_37_pe_out;
  wire       [7:0]    pE_37_acout;
  wire       [7:0]    pE_37_bcout;
  wire       [31:0]   pE_38_pe_out;
  wire       [7:0]    pE_38_acout;
  wire       [7:0]    pE_38_bcout;
  wire       [31:0]   pE_39_pe_out;
  wire       [7:0]    pE_39_acout;
  wire       [7:0]    pE_39_bcout;
  wire       [31:0]   pE_40_pe_out;
  wire       [7:0]    pE_40_acout;
  wire       [7:0]    pE_40_bcout;
  wire       [31:0]   pE_41_pe_out;
  wire       [7:0]    pE_41_acout;
  wire       [7:0]    pE_41_bcout;
  wire       [31:0]   pE_42_pe_out;
  wire       [7:0]    pE_42_acout;
  wire       [7:0]    pE_42_bcout;
  wire       [31:0]   pE_43_pe_out;
  wire       [7:0]    pE_43_acout;
  wire       [7:0]    pE_43_bcout;
  wire       [31:0]   pE_44_pe_out;
  wire       [7:0]    pE_44_acout;
  wire       [7:0]    pE_44_bcout;
  wire       [31:0]   pE_45_pe_out;
  wire       [7:0]    pE_45_acout;
  wire       [7:0]    pE_45_bcout;
  wire       [31:0]   pE_46_pe_out;
  wire       [7:0]    pE_46_acout;
  wire       [7:0]    pE_46_bcout;
  wire       [31:0]   pE_47_pe_out;
  wire       [7:0]    pE_47_acout;
  wire       [7:0]    pE_47_bcout;
  wire       [31:0]   pE_48_pe_out;
  wire       [7:0]    pE_48_acout;
  wire       [7:0]    pE_48_bcout;
  wire       [31:0]   pE_49_pe_out;
  wire       [7:0]    pE_49_acout;
  wire       [7:0]    pE_49_bcout;
  wire       [31:0]   pE_50_pe_out;
  wire       [7:0]    pE_50_acout;
  wire       [7:0]    pE_50_bcout;
  wire       [31:0]   pE_51_pe_out;
  wire       [7:0]    pE_51_acout;
  wire       [7:0]    pE_51_bcout;
  wire       [31:0]   pE_52_pe_out;
  wire       [7:0]    pE_52_acout;
  wire       [7:0]    pE_52_bcout;
  wire       [31:0]   pE_53_pe_out;
  wire       [7:0]    pE_53_acout;
  wire       [7:0]    pE_53_bcout;
  wire       [31:0]   pE_54_pe_out;
  wire       [7:0]    pE_54_acout;
  wire       [7:0]    pE_54_bcout;
  wire       [31:0]   pE_55_pe_out;
  wire       [7:0]    pE_55_acout;
  wire       [7:0]    pE_55_bcout;
  wire       [31:0]   pE_56_pe_out;
  wire       [7:0]    pE_56_acout;
  wire       [7:0]    pE_56_bcout;
  wire       [31:0]   pE_57_pe_out;
  wire       [7:0]    pE_57_acout;
  wire       [7:0]    pE_57_bcout;
  wire       [31:0]   pE_58_pe_out;
  wire       [7:0]    pE_58_acout;
  wire       [7:0]    pE_58_bcout;
  wire       [31:0]   pE_59_pe_out;
  wire       [7:0]    pE_59_acout;
  wire       [7:0]    pE_59_bcout;
  wire       [31:0]   pE_60_pe_out;
  wire       [7:0]    pE_60_acout;
  wire       [7:0]    pE_60_bcout;
  wire       [31:0]   pE_61_pe_out;
  wire       [7:0]    pE_61_acout;
  wire       [7:0]    pE_61_bcout;
  wire       [31:0]   pE_62_pe_out;
  wire       [7:0]    pE_62_acout;
  wire       [7:0]    pE_62_bcout;
  wire       [31:0]   pE_63_pe_out;
  wire       [7:0]    pE_63_acout;
  wire       [7:0]    pE_63_bcout;
  reg        [13:0]   CE_srl;
  reg        [13:0]   SCLR_srl;
  wire       [7:0]    ACOUT_0_0;
  wire       [7:0]    ACOUT_0_1;
  wire       [7:0]    ACOUT_0_2;
  wire       [7:0]    ACOUT_0_3;
  wire       [7:0]    ACOUT_0_4;
  wire       [7:0]    ACOUT_0_5;
  wire       [7:0]    ACOUT_0_6;
  wire       [7:0]    ACOUT_0_7;
  wire       [7:0]    ACOUT_1_0;
  wire       [7:0]    ACOUT_1_1;
  wire       [7:0]    ACOUT_1_2;
  wire       [7:0]    ACOUT_1_3;
  wire       [7:0]    ACOUT_1_4;
  wire       [7:0]    ACOUT_1_5;
  wire       [7:0]    ACOUT_1_6;
  wire       [7:0]    ACOUT_1_7;
  wire       [7:0]    ACOUT_2_0;
  wire       [7:0]    ACOUT_2_1;
  wire       [7:0]    ACOUT_2_2;
  wire       [7:0]    ACOUT_2_3;
  wire       [7:0]    ACOUT_2_4;
  wire       [7:0]    ACOUT_2_5;
  wire       [7:0]    ACOUT_2_6;
  wire       [7:0]    ACOUT_2_7;
  wire       [7:0]    ACOUT_3_0;
  wire       [7:0]    ACOUT_3_1;
  wire       [7:0]    ACOUT_3_2;
  wire       [7:0]    ACOUT_3_3;
  wire       [7:0]    ACOUT_3_4;
  wire       [7:0]    ACOUT_3_5;
  wire       [7:0]    ACOUT_3_6;
  wire       [7:0]    ACOUT_3_7;
  wire       [7:0]    ACOUT_4_0;
  wire       [7:0]    ACOUT_4_1;
  wire       [7:0]    ACOUT_4_2;
  wire       [7:0]    ACOUT_4_3;
  wire       [7:0]    ACOUT_4_4;
  wire       [7:0]    ACOUT_4_5;
  wire       [7:0]    ACOUT_4_6;
  wire       [7:0]    ACOUT_4_7;
  wire       [7:0]    ACOUT_5_0;
  wire       [7:0]    ACOUT_5_1;
  wire       [7:0]    ACOUT_5_2;
  wire       [7:0]    ACOUT_5_3;
  wire       [7:0]    ACOUT_5_4;
  wire       [7:0]    ACOUT_5_5;
  wire       [7:0]    ACOUT_5_6;
  wire       [7:0]    ACOUT_5_7;
  wire       [7:0]    ACOUT_6_0;
  wire       [7:0]    ACOUT_6_1;
  wire       [7:0]    ACOUT_6_2;
  wire       [7:0]    ACOUT_6_3;
  wire       [7:0]    ACOUT_6_4;
  wire       [7:0]    ACOUT_6_5;
  wire       [7:0]    ACOUT_6_6;
  wire       [7:0]    ACOUT_6_7;
  wire       [7:0]    ACOUT_7_0;
  wire       [7:0]    ACOUT_7_1;
  wire       [7:0]    ACOUT_7_2;
  wire       [7:0]    ACOUT_7_3;
  wire       [7:0]    ACOUT_7_4;
  wire       [7:0]    ACOUT_7_5;
  wire       [7:0]    ACOUT_7_6;
  wire       [7:0]    ACOUT_7_7;
  wire       [7:0]    BCOUT_0_0;
  wire       [7:0]    BCOUT_0_1;
  wire       [7:0]    BCOUT_0_2;
  wire       [7:0]    BCOUT_0_3;
  wire       [7:0]    BCOUT_0_4;
  wire       [7:0]    BCOUT_0_5;
  wire       [7:0]    BCOUT_0_6;
  wire       [7:0]    BCOUT_0_7;
  wire       [7:0]    BCOUT_1_0;
  wire       [7:0]    BCOUT_1_1;
  wire       [7:0]    BCOUT_1_2;
  wire       [7:0]    BCOUT_1_3;
  wire       [7:0]    BCOUT_1_4;
  wire       [7:0]    BCOUT_1_5;
  wire       [7:0]    BCOUT_1_6;
  wire       [7:0]    BCOUT_1_7;
  wire       [7:0]    BCOUT_2_0;
  wire       [7:0]    BCOUT_2_1;
  wire       [7:0]    BCOUT_2_2;
  wire       [7:0]    BCOUT_2_3;
  wire       [7:0]    BCOUT_2_4;
  wire       [7:0]    BCOUT_2_5;
  wire       [7:0]    BCOUT_2_6;
  wire       [7:0]    BCOUT_2_7;
  wire       [7:0]    BCOUT_3_0;
  wire       [7:0]    BCOUT_3_1;
  wire       [7:0]    BCOUT_3_2;
  wire       [7:0]    BCOUT_3_3;
  wire       [7:0]    BCOUT_3_4;
  wire       [7:0]    BCOUT_3_5;
  wire       [7:0]    BCOUT_3_6;
  wire       [7:0]    BCOUT_3_7;
  wire       [7:0]    BCOUT_4_0;
  wire       [7:0]    BCOUT_4_1;
  wire       [7:0]    BCOUT_4_2;
  wire       [7:0]    BCOUT_4_3;
  wire       [7:0]    BCOUT_4_4;
  wire       [7:0]    BCOUT_4_5;
  wire       [7:0]    BCOUT_4_6;
  wire       [7:0]    BCOUT_4_7;
  wire       [7:0]    BCOUT_5_0;
  wire       [7:0]    BCOUT_5_1;
  wire       [7:0]    BCOUT_5_2;
  wire       [7:0]    BCOUT_5_3;
  wire       [7:0]    BCOUT_5_4;
  wire       [7:0]    BCOUT_5_5;
  wire       [7:0]    BCOUT_5_6;
  wire       [7:0]    BCOUT_5_7;
  wire       [7:0]    BCOUT_6_0;
  wire       [7:0]    BCOUT_6_1;
  wire       [7:0]    BCOUT_6_2;
  wire       [7:0]    BCOUT_6_3;
  wire       [7:0]    BCOUT_6_4;
  wire       [7:0]    BCOUT_6_5;
  wire       [7:0]    BCOUT_6_6;
  wire       [7:0]    BCOUT_6_7;
  wire       [7:0]    BCOUT_7_0;
  wire       [7:0]    BCOUT_7_1;
  wire       [7:0]    BCOUT_7_2;
  wire       [7:0]    BCOUT_7_3;
  wire       [7:0]    BCOUT_7_4;
  wire       [7:0]    BCOUT_7_5;
  wire       [7:0]    BCOUT_7_6;
  wire       [7:0]    BCOUT_7_7;

  PE pe_00 (
    .clk    (clk               ), //i
    .CE     (CE                ), //i
    .SCLR   (SCLR              ), //i
    .a      (pe_00_a[7:0]      ), //i
    .b      (pe_00_b[7:0]      ), //i
    .pe_out (pe_00_pe_out[31:0]), //o
    .acout  (pe_00_acout[7:0]  ), //o
    .bcout  (pe_00_bcout[7:0]  )  //o
  );
  PE pE_1 (
    .clk    (clk              ), //i
    .CE     (pE_1_CE          ), //i
    .SCLR   (pE_1_SCLR        ), //i
    .a      (ACOUT_0_0[7:0]   ), //i
    .b      (pE_1_b[7:0]      ), //i
    .pe_out (pE_1_pe_out[31:0]), //o
    .acout  (pE_1_acout[7:0]  ), //o
    .bcout  (pE_1_bcout[7:0]  )  //o
  );
  PE pE_2 (
    .clk    (clk              ), //i
    .CE     (pE_2_CE          ), //i
    .SCLR   (pE_2_SCLR        ), //i
    .a      (ACOUT_0_1[7:0]   ), //i
    .b      (pE_2_b[7:0]      ), //i
    .pe_out (pE_2_pe_out[31:0]), //o
    .acout  (pE_2_acout[7:0]  ), //o
    .bcout  (pE_2_bcout[7:0]  )  //o
  );
  PE pE_3 (
    .clk    (clk              ), //i
    .CE     (pE_3_CE          ), //i
    .SCLR   (pE_3_SCLR        ), //i
    .a      (ACOUT_0_2[7:0]   ), //i
    .b      (pE_3_b[7:0]      ), //i
    .pe_out (pE_3_pe_out[31:0]), //o
    .acout  (pE_3_acout[7:0]  ), //o
    .bcout  (pE_3_bcout[7:0]  )  //o
  );
  PE pE_4 (
    .clk    (clk              ), //i
    .CE     (pE_4_CE          ), //i
    .SCLR   (pE_4_SCLR        ), //i
    .a      (ACOUT_0_3[7:0]   ), //i
    .b      (pE_4_b[7:0]      ), //i
    .pe_out (pE_4_pe_out[31:0]), //o
    .acout  (pE_4_acout[7:0]  ), //o
    .bcout  (pE_4_bcout[7:0]  )  //o
  );
  PE pE_5 (
    .clk    (clk              ), //i
    .CE     (pE_5_CE          ), //i
    .SCLR   (pE_5_SCLR        ), //i
    .a      (ACOUT_0_4[7:0]   ), //i
    .b      (pE_5_b[7:0]      ), //i
    .pe_out (pE_5_pe_out[31:0]), //o
    .acout  (pE_5_acout[7:0]  ), //o
    .bcout  (pE_5_bcout[7:0]  )  //o
  );
  PE pE_6 (
    .clk    (clk              ), //i
    .CE     (pE_6_CE          ), //i
    .SCLR   (pE_6_SCLR        ), //i
    .a      (ACOUT_0_5[7:0]   ), //i
    .b      (pE_6_b[7:0]      ), //i
    .pe_out (pE_6_pe_out[31:0]), //o
    .acout  (pE_6_acout[7:0]  ), //o
    .bcout  (pE_6_bcout[7:0]  )  //o
  );
  PE pE_7 (
    .clk    (clk              ), //i
    .CE     (pE_7_CE          ), //i
    .SCLR   (pE_7_SCLR        ), //i
    .a      (ACOUT_0_6[7:0]   ), //i
    .b      (pE_7_b[7:0]      ), //i
    .pe_out (pE_7_pe_out[31:0]), //o
    .acout  (pE_7_acout[7:0]  ), //o
    .bcout  (pE_7_bcout[7:0]  )  //o
  );
  PE pE_8 (
    .clk    (clk              ), //i
    .CE     (pE_8_CE          ), //i
    .SCLR   (pE_8_SCLR        ), //i
    .a      (pE_8_a[7:0]      ), //i
    .b      (BCOUT_0_0[7:0]   ), //i
    .pe_out (pE_8_pe_out[31:0]), //o
    .acout  (pE_8_acout[7:0]  ), //o
    .bcout  (pE_8_bcout[7:0]  )  //o
  );
  PE pE_9 (
    .clk    (clk              ), //i
    .CE     (pE_9_CE          ), //i
    .SCLR   (pE_9_SCLR        ), //i
    .a      (pE_9_a[7:0]      ), //i
    .b      (BCOUT_1_0[7:0]   ), //i
    .pe_out (pE_9_pe_out[31:0]), //o
    .acout  (pE_9_acout[7:0]  ), //o
    .bcout  (pE_9_bcout[7:0]  )  //o
  );
  PE pE_10 (
    .clk    (clk               ), //i
    .CE     (pE_10_CE          ), //i
    .SCLR   (pE_10_SCLR        ), //i
    .a      (pE_10_a[7:0]      ), //i
    .b      (BCOUT_2_0[7:0]    ), //i
    .pe_out (pE_10_pe_out[31:0]), //o
    .acout  (pE_10_acout[7:0]  ), //o
    .bcout  (pE_10_bcout[7:0]  )  //o
  );
  PE pE_11 (
    .clk    (clk               ), //i
    .CE     (pE_11_CE          ), //i
    .SCLR   (pE_11_SCLR        ), //i
    .a      (pE_11_a[7:0]      ), //i
    .b      (BCOUT_3_0[7:0]    ), //i
    .pe_out (pE_11_pe_out[31:0]), //o
    .acout  (pE_11_acout[7:0]  ), //o
    .bcout  (pE_11_bcout[7:0]  )  //o
  );
  PE pE_12 (
    .clk    (clk               ), //i
    .CE     (pE_12_CE          ), //i
    .SCLR   (pE_12_SCLR        ), //i
    .a      (pE_12_a[7:0]      ), //i
    .b      (BCOUT_4_0[7:0]    ), //i
    .pe_out (pE_12_pe_out[31:0]), //o
    .acout  (pE_12_acout[7:0]  ), //o
    .bcout  (pE_12_bcout[7:0]  )  //o
  );
  PE pE_13 (
    .clk    (clk               ), //i
    .CE     (pE_13_CE          ), //i
    .SCLR   (pE_13_SCLR        ), //i
    .a      (pE_13_a[7:0]      ), //i
    .b      (BCOUT_5_0[7:0]    ), //i
    .pe_out (pE_13_pe_out[31:0]), //o
    .acout  (pE_13_acout[7:0]  ), //o
    .bcout  (pE_13_bcout[7:0]  )  //o
  );
  PE pE_14 (
    .clk    (clk               ), //i
    .CE     (pE_14_CE          ), //i
    .SCLR   (pE_14_SCLR        ), //i
    .a      (pE_14_a[7:0]      ), //i
    .b      (BCOUT_6_0[7:0]    ), //i
    .pe_out (pE_14_pe_out[31:0]), //o
    .acout  (pE_14_acout[7:0]  ), //o
    .bcout  (pE_14_bcout[7:0]  )  //o
  );
  PE pE_15 (
    .clk    (clk               ), //i
    .CE     (pE_15_CE          ), //i
    .SCLR   (pE_15_SCLR        ), //i
    .a      (ACOUT_1_0[7:0]    ), //i
    .b      (BCOUT_0_1[7:0]    ), //i
    .pe_out (pE_15_pe_out[31:0]), //o
    .acout  (pE_15_acout[7:0]  ), //o
    .bcout  (pE_15_bcout[7:0]  )  //o
  );
  PE pE_16 (
    .clk    (clk               ), //i
    .CE     (pE_16_CE          ), //i
    .SCLR   (pE_16_SCLR        ), //i
    .a      (ACOUT_1_1[7:0]    ), //i
    .b      (BCOUT_0_2[7:0]    ), //i
    .pe_out (pE_16_pe_out[31:0]), //o
    .acout  (pE_16_acout[7:0]  ), //o
    .bcout  (pE_16_bcout[7:0]  )  //o
  );
  PE pE_17 (
    .clk    (clk               ), //i
    .CE     (pE_17_CE          ), //i
    .SCLR   (pE_17_SCLR        ), //i
    .a      (ACOUT_1_2[7:0]    ), //i
    .b      (BCOUT_0_3[7:0]    ), //i
    .pe_out (pE_17_pe_out[31:0]), //o
    .acout  (pE_17_acout[7:0]  ), //o
    .bcout  (pE_17_bcout[7:0]  )  //o
  );
  PE pE_18 (
    .clk    (clk               ), //i
    .CE     (pE_18_CE          ), //i
    .SCLR   (pE_18_SCLR        ), //i
    .a      (ACOUT_1_3[7:0]    ), //i
    .b      (BCOUT_0_4[7:0]    ), //i
    .pe_out (pE_18_pe_out[31:0]), //o
    .acout  (pE_18_acout[7:0]  ), //o
    .bcout  (pE_18_bcout[7:0]  )  //o
  );
  PE pE_19 (
    .clk    (clk               ), //i
    .CE     (pE_19_CE          ), //i
    .SCLR   (pE_19_SCLR        ), //i
    .a      (ACOUT_1_4[7:0]    ), //i
    .b      (BCOUT_0_5[7:0]    ), //i
    .pe_out (pE_19_pe_out[31:0]), //o
    .acout  (pE_19_acout[7:0]  ), //o
    .bcout  (pE_19_bcout[7:0]  )  //o
  );
  PE pE_20 (
    .clk    (clk               ), //i
    .CE     (pE_20_CE          ), //i
    .SCLR   (pE_20_SCLR        ), //i
    .a      (ACOUT_1_5[7:0]    ), //i
    .b      (BCOUT_0_6[7:0]    ), //i
    .pe_out (pE_20_pe_out[31:0]), //o
    .acout  (pE_20_acout[7:0]  ), //o
    .bcout  (pE_20_bcout[7:0]  )  //o
  );
  PE pE_21 (
    .clk    (clk               ), //i
    .CE     (pE_21_CE          ), //i
    .SCLR   (pE_21_SCLR        ), //i
    .a      (ACOUT_1_6[7:0]    ), //i
    .b      (BCOUT_0_7[7:0]    ), //i
    .pe_out (pE_21_pe_out[31:0]), //o
    .acout  (pE_21_acout[7:0]  ), //o
    .bcout  (pE_21_bcout[7:0]  )  //o
  );
  PE pE_22 (
    .clk    (clk               ), //i
    .CE     (pE_22_CE          ), //i
    .SCLR   (pE_22_SCLR        ), //i
    .a      (ACOUT_2_0[7:0]    ), //i
    .b      (BCOUT_1_1[7:0]    ), //i
    .pe_out (pE_22_pe_out[31:0]), //o
    .acout  (pE_22_acout[7:0]  ), //o
    .bcout  (pE_22_bcout[7:0]  )  //o
  );
  PE pE_23 (
    .clk    (clk               ), //i
    .CE     (pE_23_CE          ), //i
    .SCLR   (pE_23_SCLR        ), //i
    .a      (ACOUT_2_1[7:0]    ), //i
    .b      (BCOUT_1_2[7:0]    ), //i
    .pe_out (pE_23_pe_out[31:0]), //o
    .acout  (pE_23_acout[7:0]  ), //o
    .bcout  (pE_23_bcout[7:0]  )  //o
  );
  PE pE_24 (
    .clk    (clk               ), //i
    .CE     (pE_24_CE          ), //i
    .SCLR   (pE_24_SCLR        ), //i
    .a      (ACOUT_2_2[7:0]    ), //i
    .b      (BCOUT_1_3[7:0]    ), //i
    .pe_out (pE_24_pe_out[31:0]), //o
    .acout  (pE_24_acout[7:0]  ), //o
    .bcout  (pE_24_bcout[7:0]  )  //o
  );
  PE pE_25 (
    .clk    (clk               ), //i
    .CE     (pE_25_CE          ), //i
    .SCLR   (pE_25_SCLR        ), //i
    .a      (ACOUT_2_3[7:0]    ), //i
    .b      (BCOUT_1_4[7:0]    ), //i
    .pe_out (pE_25_pe_out[31:0]), //o
    .acout  (pE_25_acout[7:0]  ), //o
    .bcout  (pE_25_bcout[7:0]  )  //o
  );
  PE pE_26 (
    .clk    (clk               ), //i
    .CE     (pE_26_CE          ), //i
    .SCLR   (pE_26_SCLR        ), //i
    .a      (ACOUT_2_4[7:0]    ), //i
    .b      (BCOUT_1_5[7:0]    ), //i
    .pe_out (pE_26_pe_out[31:0]), //o
    .acout  (pE_26_acout[7:0]  ), //o
    .bcout  (pE_26_bcout[7:0]  )  //o
  );
  PE pE_27 (
    .clk    (clk               ), //i
    .CE     (pE_27_CE          ), //i
    .SCLR   (pE_27_SCLR        ), //i
    .a      (ACOUT_2_5[7:0]    ), //i
    .b      (BCOUT_1_6[7:0]    ), //i
    .pe_out (pE_27_pe_out[31:0]), //o
    .acout  (pE_27_acout[7:0]  ), //o
    .bcout  (pE_27_bcout[7:0]  )  //o
  );
  PE pE_28 (
    .clk    (clk               ), //i
    .CE     (pE_28_CE          ), //i
    .SCLR   (pE_28_SCLR        ), //i
    .a      (ACOUT_2_6[7:0]    ), //i
    .b      (BCOUT_1_7[7:0]    ), //i
    .pe_out (pE_28_pe_out[31:0]), //o
    .acout  (pE_28_acout[7:0]  ), //o
    .bcout  (pE_28_bcout[7:0]  )  //o
  );
  PE pE_29 (
    .clk    (clk               ), //i
    .CE     (pE_29_CE          ), //i
    .SCLR   (pE_29_SCLR        ), //i
    .a      (ACOUT_3_0[7:0]    ), //i
    .b      (BCOUT_2_1[7:0]    ), //i
    .pe_out (pE_29_pe_out[31:0]), //o
    .acout  (pE_29_acout[7:0]  ), //o
    .bcout  (pE_29_bcout[7:0]  )  //o
  );
  PE pE_30 (
    .clk    (clk               ), //i
    .CE     (pE_30_CE          ), //i
    .SCLR   (pE_30_SCLR        ), //i
    .a      (ACOUT_3_1[7:0]    ), //i
    .b      (BCOUT_2_2[7:0]    ), //i
    .pe_out (pE_30_pe_out[31:0]), //o
    .acout  (pE_30_acout[7:0]  ), //o
    .bcout  (pE_30_bcout[7:0]  )  //o
  );
  PE pE_31 (
    .clk    (clk               ), //i
    .CE     (pE_31_CE          ), //i
    .SCLR   (pE_31_SCLR        ), //i
    .a      (ACOUT_3_2[7:0]    ), //i
    .b      (BCOUT_2_3[7:0]    ), //i
    .pe_out (pE_31_pe_out[31:0]), //o
    .acout  (pE_31_acout[7:0]  ), //o
    .bcout  (pE_31_bcout[7:0]  )  //o
  );
  PE pE_32 (
    .clk    (clk               ), //i
    .CE     (pE_32_CE          ), //i
    .SCLR   (pE_32_SCLR        ), //i
    .a      (ACOUT_3_3[7:0]    ), //i
    .b      (BCOUT_2_4[7:0]    ), //i
    .pe_out (pE_32_pe_out[31:0]), //o
    .acout  (pE_32_acout[7:0]  ), //o
    .bcout  (pE_32_bcout[7:0]  )  //o
  );
  PE pE_33 (
    .clk    (clk               ), //i
    .CE     (pE_33_CE          ), //i
    .SCLR   (pE_33_SCLR        ), //i
    .a      (ACOUT_3_4[7:0]    ), //i
    .b      (BCOUT_2_5[7:0]    ), //i
    .pe_out (pE_33_pe_out[31:0]), //o
    .acout  (pE_33_acout[7:0]  ), //o
    .bcout  (pE_33_bcout[7:0]  )  //o
  );
  PE pE_34 (
    .clk    (clk               ), //i
    .CE     (pE_34_CE          ), //i
    .SCLR   (pE_34_SCLR        ), //i
    .a      (ACOUT_3_5[7:0]    ), //i
    .b      (BCOUT_2_6[7:0]    ), //i
    .pe_out (pE_34_pe_out[31:0]), //o
    .acout  (pE_34_acout[7:0]  ), //o
    .bcout  (pE_34_bcout[7:0]  )  //o
  );
  PE pE_35 (
    .clk    (clk               ), //i
    .CE     (pE_35_CE          ), //i
    .SCLR   (pE_35_SCLR        ), //i
    .a      (ACOUT_3_6[7:0]    ), //i
    .b      (BCOUT_2_7[7:0]    ), //i
    .pe_out (pE_35_pe_out[31:0]), //o
    .acout  (pE_35_acout[7:0]  ), //o
    .bcout  (pE_35_bcout[7:0]  )  //o
  );
  PE pE_36 (
    .clk    (clk               ), //i
    .CE     (pE_36_CE          ), //i
    .SCLR   (pE_36_SCLR        ), //i
    .a      (ACOUT_4_0[7:0]    ), //i
    .b      (BCOUT_3_1[7:0]    ), //i
    .pe_out (pE_36_pe_out[31:0]), //o
    .acout  (pE_36_acout[7:0]  ), //o
    .bcout  (pE_36_bcout[7:0]  )  //o
  );
  PE pE_37 (
    .clk    (clk               ), //i
    .CE     (pE_37_CE          ), //i
    .SCLR   (pE_37_SCLR        ), //i
    .a      (ACOUT_4_1[7:0]    ), //i
    .b      (BCOUT_3_2[7:0]    ), //i
    .pe_out (pE_37_pe_out[31:0]), //o
    .acout  (pE_37_acout[7:0]  ), //o
    .bcout  (pE_37_bcout[7:0]  )  //o
  );
  PE pE_38 (
    .clk    (clk               ), //i
    .CE     (pE_38_CE          ), //i
    .SCLR   (pE_38_SCLR        ), //i
    .a      (ACOUT_4_2[7:0]    ), //i
    .b      (BCOUT_3_3[7:0]    ), //i
    .pe_out (pE_38_pe_out[31:0]), //o
    .acout  (pE_38_acout[7:0]  ), //o
    .bcout  (pE_38_bcout[7:0]  )  //o
  );
  PE pE_39 (
    .clk    (clk               ), //i
    .CE     (pE_39_CE          ), //i
    .SCLR   (pE_39_SCLR        ), //i
    .a      (ACOUT_4_3[7:0]    ), //i
    .b      (BCOUT_3_4[7:0]    ), //i
    .pe_out (pE_39_pe_out[31:0]), //o
    .acout  (pE_39_acout[7:0]  ), //o
    .bcout  (pE_39_bcout[7:0]  )  //o
  );
  PE pE_40 (
    .clk    (clk               ), //i
    .CE     (pE_40_CE          ), //i
    .SCLR   (pE_40_SCLR        ), //i
    .a      (ACOUT_4_4[7:0]    ), //i
    .b      (BCOUT_3_5[7:0]    ), //i
    .pe_out (pE_40_pe_out[31:0]), //o
    .acout  (pE_40_acout[7:0]  ), //o
    .bcout  (pE_40_bcout[7:0]  )  //o
  );
  PE pE_41 (
    .clk    (clk               ), //i
    .CE     (pE_41_CE          ), //i
    .SCLR   (pE_41_SCLR        ), //i
    .a      (ACOUT_4_5[7:0]    ), //i
    .b      (BCOUT_3_6[7:0]    ), //i
    .pe_out (pE_41_pe_out[31:0]), //o
    .acout  (pE_41_acout[7:0]  ), //o
    .bcout  (pE_41_bcout[7:0]  )  //o
  );
  PE pE_42 (
    .clk    (clk               ), //i
    .CE     (pE_42_CE          ), //i
    .SCLR   (pE_42_SCLR        ), //i
    .a      (ACOUT_4_6[7:0]    ), //i
    .b      (BCOUT_3_7[7:0]    ), //i
    .pe_out (pE_42_pe_out[31:0]), //o
    .acout  (pE_42_acout[7:0]  ), //o
    .bcout  (pE_42_bcout[7:0]  )  //o
  );
  PE pE_43 (
    .clk    (clk               ), //i
    .CE     (pE_43_CE          ), //i
    .SCLR   (pE_43_SCLR        ), //i
    .a      (ACOUT_5_0[7:0]    ), //i
    .b      (BCOUT_4_1[7:0]    ), //i
    .pe_out (pE_43_pe_out[31:0]), //o
    .acout  (pE_43_acout[7:0]  ), //o
    .bcout  (pE_43_bcout[7:0]  )  //o
  );
  PE pE_44 (
    .clk    (clk               ), //i
    .CE     (pE_44_CE          ), //i
    .SCLR   (pE_44_SCLR        ), //i
    .a      (ACOUT_5_1[7:0]    ), //i
    .b      (BCOUT_4_2[7:0]    ), //i
    .pe_out (pE_44_pe_out[31:0]), //o
    .acout  (pE_44_acout[7:0]  ), //o
    .bcout  (pE_44_bcout[7:0]  )  //o
  );
  PE pE_45 (
    .clk    (clk               ), //i
    .CE     (pE_45_CE          ), //i
    .SCLR   (pE_45_SCLR        ), //i
    .a      (ACOUT_5_2[7:0]    ), //i
    .b      (BCOUT_4_3[7:0]    ), //i
    .pe_out (pE_45_pe_out[31:0]), //o
    .acout  (pE_45_acout[7:0]  ), //o
    .bcout  (pE_45_bcout[7:0]  )  //o
  );
  PE pE_46 (
    .clk    (clk               ), //i
    .CE     (pE_46_CE          ), //i
    .SCLR   (pE_46_SCLR        ), //i
    .a      (ACOUT_5_3[7:0]    ), //i
    .b      (BCOUT_4_4[7:0]    ), //i
    .pe_out (pE_46_pe_out[31:0]), //o
    .acout  (pE_46_acout[7:0]  ), //o
    .bcout  (pE_46_bcout[7:0]  )  //o
  );
  PE pE_47 (
    .clk    (clk               ), //i
    .CE     (pE_47_CE          ), //i
    .SCLR   (pE_47_SCLR        ), //i
    .a      (ACOUT_5_4[7:0]    ), //i
    .b      (BCOUT_4_5[7:0]    ), //i
    .pe_out (pE_47_pe_out[31:0]), //o
    .acout  (pE_47_acout[7:0]  ), //o
    .bcout  (pE_47_bcout[7:0]  )  //o
  );
  PE pE_48 (
    .clk    (clk               ), //i
    .CE     (pE_48_CE          ), //i
    .SCLR   (pE_48_SCLR        ), //i
    .a      (ACOUT_5_5[7:0]    ), //i
    .b      (BCOUT_4_6[7:0]    ), //i
    .pe_out (pE_48_pe_out[31:0]), //o
    .acout  (pE_48_acout[7:0]  ), //o
    .bcout  (pE_48_bcout[7:0]  )  //o
  );
  PE pE_49 (
    .clk    (clk               ), //i
    .CE     (pE_49_CE          ), //i
    .SCLR   (pE_49_SCLR        ), //i
    .a      (ACOUT_5_6[7:0]    ), //i
    .b      (BCOUT_4_7[7:0]    ), //i
    .pe_out (pE_49_pe_out[31:0]), //o
    .acout  (pE_49_acout[7:0]  ), //o
    .bcout  (pE_49_bcout[7:0]  )  //o
  );
  PE pE_50 (
    .clk    (clk               ), //i
    .CE     (pE_50_CE          ), //i
    .SCLR   (pE_50_SCLR        ), //i
    .a      (ACOUT_6_0[7:0]    ), //i
    .b      (BCOUT_5_1[7:0]    ), //i
    .pe_out (pE_50_pe_out[31:0]), //o
    .acout  (pE_50_acout[7:0]  ), //o
    .bcout  (pE_50_bcout[7:0]  )  //o
  );
  PE pE_51 (
    .clk    (clk               ), //i
    .CE     (pE_51_CE          ), //i
    .SCLR   (pE_51_SCLR        ), //i
    .a      (ACOUT_6_1[7:0]    ), //i
    .b      (BCOUT_5_2[7:0]    ), //i
    .pe_out (pE_51_pe_out[31:0]), //o
    .acout  (pE_51_acout[7:0]  ), //o
    .bcout  (pE_51_bcout[7:0]  )  //o
  );
  PE pE_52 (
    .clk    (clk               ), //i
    .CE     (pE_52_CE          ), //i
    .SCLR   (pE_52_SCLR        ), //i
    .a      (ACOUT_6_2[7:0]    ), //i
    .b      (BCOUT_5_3[7:0]    ), //i
    .pe_out (pE_52_pe_out[31:0]), //o
    .acout  (pE_52_acout[7:0]  ), //o
    .bcout  (pE_52_bcout[7:0]  )  //o
  );
  PE pE_53 (
    .clk    (clk               ), //i
    .CE     (pE_53_CE          ), //i
    .SCLR   (pE_53_SCLR        ), //i
    .a      (ACOUT_6_3[7:0]    ), //i
    .b      (BCOUT_5_4[7:0]    ), //i
    .pe_out (pE_53_pe_out[31:0]), //o
    .acout  (pE_53_acout[7:0]  ), //o
    .bcout  (pE_53_bcout[7:0]  )  //o
  );
  PE pE_54 (
    .clk    (clk               ), //i
    .CE     (pE_54_CE          ), //i
    .SCLR   (pE_54_SCLR        ), //i
    .a      (ACOUT_6_4[7:0]    ), //i
    .b      (BCOUT_5_5[7:0]    ), //i
    .pe_out (pE_54_pe_out[31:0]), //o
    .acout  (pE_54_acout[7:0]  ), //o
    .bcout  (pE_54_bcout[7:0]  )  //o
  );
  PE pE_55 (
    .clk    (clk               ), //i
    .CE     (pE_55_CE          ), //i
    .SCLR   (pE_55_SCLR        ), //i
    .a      (ACOUT_6_5[7:0]    ), //i
    .b      (BCOUT_5_6[7:0]    ), //i
    .pe_out (pE_55_pe_out[31:0]), //o
    .acout  (pE_55_acout[7:0]  ), //o
    .bcout  (pE_55_bcout[7:0]  )  //o
  );
  PE pE_56 (
    .clk    (clk               ), //i
    .CE     (pE_56_CE          ), //i
    .SCLR   (pE_56_SCLR        ), //i
    .a      (ACOUT_6_6[7:0]    ), //i
    .b      (BCOUT_5_7[7:0]    ), //i
    .pe_out (pE_56_pe_out[31:0]), //o
    .acout  (pE_56_acout[7:0]  ), //o
    .bcout  (pE_56_bcout[7:0]  )  //o
  );
  PE pE_57 (
    .clk    (clk               ), //i
    .CE     (pE_57_CE          ), //i
    .SCLR   (pE_57_SCLR        ), //i
    .a      (ACOUT_7_0[7:0]    ), //i
    .b      (BCOUT_6_1[7:0]    ), //i
    .pe_out (pE_57_pe_out[31:0]), //o
    .acout  (pE_57_acout[7:0]  ), //o
    .bcout  (pE_57_bcout[7:0]  )  //o
  );
  PE pE_58 (
    .clk    (clk               ), //i
    .CE     (pE_58_CE          ), //i
    .SCLR   (pE_58_SCLR        ), //i
    .a      (ACOUT_7_1[7:0]    ), //i
    .b      (BCOUT_6_2[7:0]    ), //i
    .pe_out (pE_58_pe_out[31:0]), //o
    .acout  (pE_58_acout[7:0]  ), //o
    .bcout  (pE_58_bcout[7:0]  )  //o
  );
  PE pE_59 (
    .clk    (clk               ), //i
    .CE     (pE_59_CE          ), //i
    .SCLR   (pE_59_SCLR        ), //i
    .a      (ACOUT_7_2[7:0]    ), //i
    .b      (BCOUT_6_3[7:0]    ), //i
    .pe_out (pE_59_pe_out[31:0]), //o
    .acout  (pE_59_acout[7:0]  ), //o
    .bcout  (pE_59_bcout[7:0]  )  //o
  );
  PE pE_60 (
    .clk    (clk               ), //i
    .CE     (pE_60_CE          ), //i
    .SCLR   (pE_60_SCLR        ), //i
    .a      (ACOUT_7_3[7:0]    ), //i
    .b      (BCOUT_6_4[7:0]    ), //i
    .pe_out (pE_60_pe_out[31:0]), //o
    .acout  (pE_60_acout[7:0]  ), //o
    .bcout  (pE_60_bcout[7:0]  )  //o
  );
  PE pE_61 (
    .clk    (clk               ), //i
    .CE     (pE_61_CE          ), //i
    .SCLR   (pE_61_SCLR        ), //i
    .a      (ACOUT_7_4[7:0]    ), //i
    .b      (BCOUT_6_5[7:0]    ), //i
    .pe_out (pE_61_pe_out[31:0]), //o
    .acout  (pE_61_acout[7:0]  ), //o
    .bcout  (pE_61_bcout[7:0]  )  //o
  );
  PE pE_62 (
    .clk    (clk               ), //i
    .CE     (pE_62_CE          ), //i
    .SCLR   (pE_62_SCLR        ), //i
    .a      (ACOUT_7_5[7:0]    ), //i
    .b      (BCOUT_6_6[7:0]    ), //i
    .pe_out (pE_62_pe_out[31:0]), //o
    .acout  (pE_62_acout[7:0]  ), //o
    .bcout  (pE_62_bcout[7:0]  )  //o
  );
  PE pE_63 (
    .clk    (clk               ), //i
    .CE     (pE_63_CE          ), //i
    .SCLR   (pE_63_SCLR        ), //i
    .a      (ACOUT_7_6[7:0]    ), //i
    .b      (BCOUT_6_7[7:0]    ), //i
    .pe_out (pE_63_pe_out[31:0]), //o
    .acout  (pE_63_acout[7:0]  ), //o
    .bcout  (pE_63_bcout[7:0]  )  //o
  );
  assign pe_00_a = A[7 : 0];
  assign pe_00_b = B[7 : 0];
  always @(*) begin
    Tile_OUT[31 : 0] = pe_00_pe_out;
    Tile_OUT[63 : 32] = pE_1_pe_out;
    Tile_OUT[95 : 64] = pE_2_pe_out;
    Tile_OUT[127 : 96] = pE_3_pe_out;
    Tile_OUT[159 : 128] = pE_4_pe_out;
    Tile_OUT[191 : 160] = pE_5_pe_out;
    Tile_OUT[223 : 192] = pE_6_pe_out;
    Tile_OUT[255 : 224] = pE_7_pe_out;
    Tile_OUT[287 : 256] = pE_8_pe_out;
    Tile_OUT[543 : 512] = pE_9_pe_out;
    Tile_OUT[799 : 768] = pE_10_pe_out;
    Tile_OUT[1055 : 1024] = pE_11_pe_out;
    Tile_OUT[1311 : 1280] = pE_12_pe_out;
    Tile_OUT[1567 : 1536] = pE_13_pe_out;
    Tile_OUT[1823 : 1792] = pE_14_pe_out;
    Tile_OUT[319 : 288] = pE_15_pe_out;
    Tile_OUT[575 : 544] = pE_16_pe_out;
    Tile_OUT[831 : 800] = pE_17_pe_out;
    Tile_OUT[1087 : 1056] = pE_18_pe_out;
    Tile_OUT[1343 : 1312] = pE_19_pe_out;
    Tile_OUT[1599 : 1568] = pE_20_pe_out;
    Tile_OUT[1855 : 1824] = pE_21_pe_out;
    Tile_OUT[351 : 320] = pE_22_pe_out;
    Tile_OUT[607 : 576] = pE_23_pe_out;
    Tile_OUT[863 : 832] = pE_24_pe_out;
    Tile_OUT[1119 : 1088] = pE_25_pe_out;
    Tile_OUT[1375 : 1344] = pE_26_pe_out;
    Tile_OUT[1631 : 1600] = pE_27_pe_out;
    Tile_OUT[1887 : 1856] = pE_28_pe_out;
    Tile_OUT[383 : 352] = pE_29_pe_out;
    Tile_OUT[639 : 608] = pE_30_pe_out;
    Tile_OUT[895 : 864] = pE_31_pe_out;
    Tile_OUT[1151 : 1120] = pE_32_pe_out;
    Tile_OUT[1407 : 1376] = pE_33_pe_out;
    Tile_OUT[1663 : 1632] = pE_34_pe_out;
    Tile_OUT[1919 : 1888] = pE_35_pe_out;
    Tile_OUT[415 : 384] = pE_36_pe_out;
    Tile_OUT[671 : 640] = pE_37_pe_out;
    Tile_OUT[927 : 896] = pE_38_pe_out;
    Tile_OUT[1183 : 1152] = pE_39_pe_out;
    Tile_OUT[1439 : 1408] = pE_40_pe_out;
    Tile_OUT[1695 : 1664] = pE_41_pe_out;
    Tile_OUT[1951 : 1920] = pE_42_pe_out;
    Tile_OUT[447 : 416] = pE_43_pe_out;
    Tile_OUT[703 : 672] = pE_44_pe_out;
    Tile_OUT[959 : 928] = pE_45_pe_out;
    Tile_OUT[1215 : 1184] = pE_46_pe_out;
    Tile_OUT[1471 : 1440] = pE_47_pe_out;
    Tile_OUT[1727 : 1696] = pE_48_pe_out;
    Tile_OUT[1983 : 1952] = pE_49_pe_out;
    Tile_OUT[479 : 448] = pE_50_pe_out;
    Tile_OUT[735 : 704] = pE_51_pe_out;
    Tile_OUT[991 : 960] = pE_52_pe_out;
    Tile_OUT[1247 : 1216] = pE_53_pe_out;
    Tile_OUT[1503 : 1472] = pE_54_pe_out;
    Tile_OUT[1759 : 1728] = pE_55_pe_out;
    Tile_OUT[2015 : 1984] = pE_56_pe_out;
    Tile_OUT[511 : 480] = pE_57_pe_out;
    Tile_OUT[767 : 736] = pE_58_pe_out;
    Tile_OUT[1023 : 992] = pE_59_pe_out;
    Tile_OUT[1279 : 1248] = pE_60_pe_out;
    Tile_OUT[1535 : 1504] = pE_61_pe_out;
    Tile_OUT[1791 : 1760] = pE_62_pe_out;
    Tile_OUT[2047 : 2016] = pE_63_pe_out;
  end

  assign ACOUT_0_0 = pe_00_acout;
  assign BCOUT_0_0 = pe_00_bcout;
  assign pE_1_CE = CE_srl[0];
  assign pE_1_SCLR = SCLR_srl[0];
  assign pE_1_b = B[15 : 8];
  assign ACOUT_0_1 = pE_1_acout;
  assign BCOUT_0_1 = pE_1_bcout;
  assign pE_2_CE = CE_srl[1];
  assign pE_2_SCLR = SCLR_srl[1];
  assign pE_2_b = B[23 : 16];
  assign ACOUT_0_2 = pE_2_acout;
  assign BCOUT_0_2 = pE_2_bcout;
  assign pE_3_CE = CE_srl[2];
  assign pE_3_SCLR = SCLR_srl[2];
  assign pE_3_b = B[31 : 24];
  assign ACOUT_0_3 = pE_3_acout;
  assign BCOUT_0_3 = pE_3_bcout;
  assign pE_4_CE = CE_srl[3];
  assign pE_4_SCLR = SCLR_srl[3];
  assign pE_4_b = B[39 : 32];
  assign ACOUT_0_4 = pE_4_acout;
  assign BCOUT_0_4 = pE_4_bcout;
  assign pE_5_CE = CE_srl[4];
  assign pE_5_SCLR = SCLR_srl[4];
  assign pE_5_b = B[47 : 40];
  assign ACOUT_0_5 = pE_5_acout;
  assign BCOUT_0_5 = pE_5_bcout;
  assign pE_6_CE = CE_srl[5];
  assign pE_6_SCLR = SCLR_srl[5];
  assign pE_6_b = B[55 : 48];
  assign ACOUT_0_6 = pE_6_acout;
  assign BCOUT_0_6 = pE_6_bcout;
  assign pE_7_CE = CE_srl[6];
  assign pE_7_SCLR = SCLR_srl[6];
  assign pE_7_b = B[63 : 56];
  assign ACOUT_0_7 = pE_7_acout;
  assign BCOUT_0_7 = pE_7_bcout;
  assign pE_8_CE = CE_srl[0];
  assign pE_8_SCLR = SCLR_srl[0];
  assign pE_8_a = A[15 : 8];
  assign ACOUT_1_0 = pE_8_acout;
  assign BCOUT_1_0 = pE_8_bcout;
  assign pE_9_CE = CE_srl[1];
  assign pE_9_SCLR = SCLR_srl[1];
  assign pE_9_a = A[23 : 16];
  assign ACOUT_2_0 = pE_9_acout;
  assign BCOUT_2_0 = pE_9_bcout;
  assign pE_10_CE = CE_srl[2];
  assign pE_10_SCLR = SCLR_srl[2];
  assign pE_10_a = A[31 : 24];
  assign ACOUT_3_0 = pE_10_acout;
  assign BCOUT_3_0 = pE_10_bcout;
  assign pE_11_CE = CE_srl[3];
  assign pE_11_SCLR = SCLR_srl[3];
  assign pE_11_a = A[39 : 32];
  assign ACOUT_4_0 = pE_11_acout;
  assign BCOUT_4_0 = pE_11_bcout;
  assign pE_12_CE = CE_srl[4];
  assign pE_12_SCLR = SCLR_srl[4];
  assign pE_12_a = A[47 : 40];
  assign ACOUT_5_0 = pE_12_acout;
  assign BCOUT_5_0 = pE_12_bcout;
  assign pE_13_CE = CE_srl[5];
  assign pE_13_SCLR = SCLR_srl[5];
  assign pE_13_a = A[55 : 48];
  assign ACOUT_6_0 = pE_13_acout;
  assign BCOUT_6_0 = pE_13_bcout;
  assign pE_14_CE = CE_srl[6];
  assign pE_14_SCLR = SCLR_srl[6];
  assign pE_14_a = A[63 : 56];
  assign ACOUT_7_0 = pE_14_acout;
  assign BCOUT_7_0 = pE_14_bcout;
  assign pE_15_CE = CE_srl[1];
  assign pE_15_SCLR = SCLR_srl[1];
  assign ACOUT_1_1 = pE_15_acout;
  assign BCOUT_1_1 = pE_15_bcout;
  assign pE_16_CE = CE_srl[2];
  assign pE_16_SCLR = SCLR_srl[2];
  assign ACOUT_1_2 = pE_16_acout;
  assign BCOUT_1_2 = pE_16_bcout;
  assign pE_17_CE = CE_srl[3];
  assign pE_17_SCLR = SCLR_srl[3];
  assign ACOUT_1_3 = pE_17_acout;
  assign BCOUT_1_3 = pE_17_bcout;
  assign pE_18_CE = CE_srl[4];
  assign pE_18_SCLR = SCLR_srl[4];
  assign ACOUT_1_4 = pE_18_acout;
  assign BCOUT_1_4 = pE_18_bcout;
  assign pE_19_CE = CE_srl[5];
  assign pE_19_SCLR = SCLR_srl[5];
  assign ACOUT_1_5 = pE_19_acout;
  assign BCOUT_1_5 = pE_19_bcout;
  assign pE_20_CE = CE_srl[6];
  assign pE_20_SCLR = SCLR_srl[6];
  assign ACOUT_1_6 = pE_20_acout;
  assign BCOUT_1_6 = pE_20_bcout;
  assign pE_21_CE = CE_srl[7];
  assign pE_21_SCLR = SCLR_srl[7];
  assign ACOUT_1_7 = pE_21_acout;
  assign BCOUT_1_7 = pE_21_bcout;
  assign pE_22_CE = CE_srl[2];
  assign pE_22_SCLR = SCLR_srl[2];
  assign ACOUT_2_1 = pE_22_acout;
  assign BCOUT_2_1 = pE_22_bcout;
  assign pE_23_CE = CE_srl[3];
  assign pE_23_SCLR = SCLR_srl[3];
  assign ACOUT_2_2 = pE_23_acout;
  assign BCOUT_2_2 = pE_23_bcout;
  assign pE_24_CE = CE_srl[4];
  assign pE_24_SCLR = SCLR_srl[4];
  assign ACOUT_2_3 = pE_24_acout;
  assign BCOUT_2_3 = pE_24_bcout;
  assign pE_25_CE = CE_srl[5];
  assign pE_25_SCLR = SCLR_srl[5];
  assign ACOUT_2_4 = pE_25_acout;
  assign BCOUT_2_4 = pE_25_bcout;
  assign pE_26_CE = CE_srl[6];
  assign pE_26_SCLR = SCLR_srl[6];
  assign ACOUT_2_5 = pE_26_acout;
  assign BCOUT_2_5 = pE_26_bcout;
  assign pE_27_CE = CE_srl[7];
  assign pE_27_SCLR = SCLR_srl[7];
  assign ACOUT_2_6 = pE_27_acout;
  assign BCOUT_2_6 = pE_27_bcout;
  assign pE_28_CE = CE_srl[8];
  assign pE_28_SCLR = SCLR_srl[8];
  assign ACOUT_2_7 = pE_28_acout;
  assign BCOUT_2_7 = pE_28_bcout;
  assign pE_29_CE = CE_srl[3];
  assign pE_29_SCLR = SCLR_srl[3];
  assign ACOUT_3_1 = pE_29_acout;
  assign BCOUT_3_1 = pE_29_bcout;
  assign pE_30_CE = CE_srl[4];
  assign pE_30_SCLR = SCLR_srl[4];
  assign ACOUT_3_2 = pE_30_acout;
  assign BCOUT_3_2 = pE_30_bcout;
  assign pE_31_CE = CE_srl[5];
  assign pE_31_SCLR = SCLR_srl[5];
  assign ACOUT_3_3 = pE_31_acout;
  assign BCOUT_3_3 = pE_31_bcout;
  assign pE_32_CE = CE_srl[6];
  assign pE_32_SCLR = SCLR_srl[6];
  assign ACOUT_3_4 = pE_32_acout;
  assign BCOUT_3_4 = pE_32_bcout;
  assign pE_33_CE = CE_srl[7];
  assign pE_33_SCLR = SCLR_srl[7];
  assign ACOUT_3_5 = pE_33_acout;
  assign BCOUT_3_5 = pE_33_bcout;
  assign pE_34_CE = CE_srl[8];
  assign pE_34_SCLR = SCLR_srl[8];
  assign ACOUT_3_6 = pE_34_acout;
  assign BCOUT_3_6 = pE_34_bcout;
  assign pE_35_CE = CE_srl[9];
  assign pE_35_SCLR = SCLR_srl[9];
  assign ACOUT_3_7 = pE_35_acout;
  assign BCOUT_3_7 = pE_35_bcout;
  assign pE_36_CE = CE_srl[4];
  assign pE_36_SCLR = SCLR_srl[4];
  assign ACOUT_4_1 = pE_36_acout;
  assign BCOUT_4_1 = pE_36_bcout;
  assign pE_37_CE = CE_srl[5];
  assign pE_37_SCLR = SCLR_srl[5];
  assign ACOUT_4_2 = pE_37_acout;
  assign BCOUT_4_2 = pE_37_bcout;
  assign pE_38_CE = CE_srl[6];
  assign pE_38_SCLR = SCLR_srl[6];
  assign ACOUT_4_3 = pE_38_acout;
  assign BCOUT_4_3 = pE_38_bcout;
  assign pE_39_CE = CE_srl[7];
  assign pE_39_SCLR = SCLR_srl[7];
  assign ACOUT_4_4 = pE_39_acout;
  assign BCOUT_4_4 = pE_39_bcout;
  assign pE_40_CE = CE_srl[8];
  assign pE_40_SCLR = SCLR_srl[8];
  assign ACOUT_4_5 = pE_40_acout;
  assign BCOUT_4_5 = pE_40_bcout;
  assign pE_41_CE = CE_srl[9];
  assign pE_41_SCLR = SCLR_srl[9];
  assign ACOUT_4_6 = pE_41_acout;
  assign BCOUT_4_6 = pE_41_bcout;
  assign pE_42_CE = CE_srl[10];
  assign pE_42_SCLR = SCLR_srl[10];
  assign ACOUT_4_7 = pE_42_acout;
  assign BCOUT_4_7 = pE_42_bcout;
  assign pE_43_CE = CE_srl[5];
  assign pE_43_SCLR = SCLR_srl[5];
  assign ACOUT_5_1 = pE_43_acout;
  assign BCOUT_5_1 = pE_43_bcout;
  assign pE_44_CE = CE_srl[6];
  assign pE_44_SCLR = SCLR_srl[6];
  assign ACOUT_5_2 = pE_44_acout;
  assign BCOUT_5_2 = pE_44_bcout;
  assign pE_45_CE = CE_srl[7];
  assign pE_45_SCLR = SCLR_srl[7];
  assign ACOUT_5_3 = pE_45_acout;
  assign BCOUT_5_3 = pE_45_bcout;
  assign pE_46_CE = CE_srl[8];
  assign pE_46_SCLR = SCLR_srl[8];
  assign ACOUT_5_4 = pE_46_acout;
  assign BCOUT_5_4 = pE_46_bcout;
  assign pE_47_CE = CE_srl[9];
  assign pE_47_SCLR = SCLR_srl[9];
  assign ACOUT_5_5 = pE_47_acout;
  assign BCOUT_5_5 = pE_47_bcout;
  assign pE_48_CE = CE_srl[10];
  assign pE_48_SCLR = SCLR_srl[10];
  assign ACOUT_5_6 = pE_48_acout;
  assign BCOUT_5_6 = pE_48_bcout;
  assign pE_49_CE = CE_srl[11];
  assign pE_49_SCLR = SCLR_srl[11];
  assign ACOUT_5_7 = pE_49_acout;
  assign BCOUT_5_7 = pE_49_bcout;
  assign pE_50_CE = CE_srl[6];
  assign pE_50_SCLR = SCLR_srl[6];
  assign ACOUT_6_1 = pE_50_acout;
  assign BCOUT_6_1 = pE_50_bcout;
  assign pE_51_CE = CE_srl[7];
  assign pE_51_SCLR = SCLR_srl[7];
  assign ACOUT_6_2 = pE_51_acout;
  assign BCOUT_6_2 = pE_51_bcout;
  assign pE_52_CE = CE_srl[8];
  assign pE_52_SCLR = SCLR_srl[8];
  assign ACOUT_6_3 = pE_52_acout;
  assign BCOUT_6_3 = pE_52_bcout;
  assign pE_53_CE = CE_srl[9];
  assign pE_53_SCLR = SCLR_srl[9];
  assign ACOUT_6_4 = pE_53_acout;
  assign BCOUT_6_4 = pE_53_bcout;
  assign pE_54_CE = CE_srl[10];
  assign pE_54_SCLR = SCLR_srl[10];
  assign ACOUT_6_5 = pE_54_acout;
  assign BCOUT_6_5 = pE_54_bcout;
  assign pE_55_CE = CE_srl[11];
  assign pE_55_SCLR = SCLR_srl[11];
  assign ACOUT_6_6 = pE_55_acout;
  assign BCOUT_6_6 = pE_55_bcout;
  assign pE_56_CE = CE_srl[12];
  assign pE_56_SCLR = SCLR_srl[12];
  assign ACOUT_6_7 = pE_56_acout;
  assign BCOUT_6_7 = pE_56_bcout;
  assign pE_57_CE = CE_srl[7];
  assign pE_57_SCLR = SCLR_srl[7];
  assign ACOUT_7_1 = pE_57_acout;
  assign BCOUT_7_1 = pE_57_bcout;
  assign pE_58_CE = CE_srl[8];
  assign pE_58_SCLR = SCLR_srl[8];
  assign ACOUT_7_2 = pE_58_acout;
  assign BCOUT_7_2 = pE_58_bcout;
  assign pE_59_CE = CE_srl[9];
  assign pE_59_SCLR = SCLR_srl[9];
  assign ACOUT_7_3 = pE_59_acout;
  assign BCOUT_7_3 = pE_59_bcout;
  assign pE_60_CE = CE_srl[10];
  assign pE_60_SCLR = SCLR_srl[10];
  assign ACOUT_7_4 = pE_60_acout;
  assign BCOUT_7_4 = pE_60_bcout;
  assign pE_61_CE = CE_srl[11];
  assign pE_61_SCLR = SCLR_srl[11];
  assign ACOUT_7_5 = pE_61_acout;
  assign BCOUT_7_5 = pE_61_bcout;
  assign pE_62_CE = CE_srl[12];
  assign pE_62_SCLR = SCLR_srl[12];
  assign ACOUT_7_6 = pE_62_acout;
  assign BCOUT_7_6 = pE_62_bcout;
  assign pE_63_CE = CE_srl[13];
  assign pE_63_SCLR = SCLR_srl[13];
  assign ACOUT_7_7 = pE_63_acout;
  assign BCOUT_7_7 = pE_63_bcout;
  always @(posedge clk) begin
    if(reset) begin
      CE_srl <= 14'h0;
      SCLR_srl <= 14'h0;
    end else begin
      CE_srl[0] <= CE;
      CE_srl[1] <= CE_srl[0];
      CE_srl[2] <= CE_srl[1];
      CE_srl[3] <= CE_srl[2];
      CE_srl[4] <= CE_srl[3];
      CE_srl[5] <= CE_srl[4];
      CE_srl[6] <= CE_srl[5];
      CE_srl[7] <= CE_srl[6];
      CE_srl[8] <= CE_srl[7];
      CE_srl[9] <= CE_srl[8];
      CE_srl[10] <= CE_srl[9];
      CE_srl[11] <= CE_srl[10];
      CE_srl[12] <= CE_srl[11];
      CE_srl[13] <= CE_srl[12];
      SCLR_srl[0] <= SCLR;
      SCLR_srl[1] <= SCLR_srl[0];
      SCLR_srl[2] <= SCLR_srl[1];
      SCLR_srl[3] <= SCLR_srl[2];
      SCLR_srl[4] <= SCLR_srl[3];
      SCLR_srl[5] <= SCLR_srl[4];
      SCLR_srl[6] <= SCLR_srl[5];
      SCLR_srl[7] <= SCLR_srl[6];
      SCLR_srl[8] <= SCLR_srl[7];
      SCLR_srl[9] <= SCLR_srl[8];
      SCLR_srl[10] <= SCLR_srl[9];
      SCLR_srl[11] <= SCLR_srl[10];
      SCLR_srl[12] <= SCLR_srl[11];
      SCLR_srl[13] <= SCLR_srl[12];
    end
  end


endmodule

module PE(
        	input clk,
        	input	CE,
        	input SCLR,
        	input	[7:0]	a,
        	input	[7:0]	b,
        	output	[31:0]	pe_out,
        	output	 [7:0]	acout,
        	output   [7:0]	bcout
        );
	    wire signed	[7:0]	a_in;
	    assign a_in = $signed(a);
          pe pe_u (
            .CLK(clk),      // input wire CLK
            .CE(CE),        // input wire CE
            .A(a_in),          // input wire [7 : 0] A
            .B({1'b0,b}),          // input wire [8 : 0] B
            .ACOUT(acout),  // output wire [29 : 0] ACOUT
            .BCOUT(bcout),  // output wire [17 : 0] BCOUT
            .P(pe_out),          // output wire [47 : 0] P
            .SCLR(SCLR)  // input wire SCLRP
	        );

endmodule
      
